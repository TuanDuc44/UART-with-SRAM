magic
tech sky130A
timestamp 1745938526
<< viali >>
rect 15948 29792 15965 29809
rect 15999 29690 16016 29707
rect 10272 29554 10289 29571
rect 11698 29554 11715 29571
rect 15700 29554 15717 29571
rect 16114 29520 16131 29537
rect 16252 29520 16269 29537
rect 10272 29486 10289 29503
rect 10410 29486 10427 29503
rect 11836 29486 11853 29503
rect 12066 29486 12083 29503
rect 12158 29486 12175 29503
rect 15792 29486 15809 29503
rect 15838 29486 15855 29503
rect 16160 29486 16177 29503
rect 11698 29452 11715 29469
rect 15700 29452 15717 29469
rect 10364 29418 10381 29435
rect 11790 29418 11807 29435
rect 12112 29418 12129 29435
rect 15792 29418 15809 29435
rect 16252 29418 16269 29435
rect 14596 29316 14613 29333
rect 15700 29316 15717 29333
rect 16620 29316 16637 29333
rect 7033 29282 7050 29299
rect 10130 29282 10147 29299
rect 11786 29282 11803 29299
rect 15144 29282 15161 29299
rect 6977 29248 6994 29265
rect 8892 29248 8909 29265
rect 8984 29248 9001 29265
rect 9996 29248 10013 29265
rect 11652 29248 11669 29265
rect 13304 29248 13321 29265
rect 14550 29248 14567 29265
rect 14734 29248 14751 29265
rect 16064 29248 16081 29265
rect 6822 29214 6839 29231
rect 13170 29214 13187 29231
rect 14642 29214 14659 29231
rect 15010 29214 15027 29231
rect 15930 29214 15947 29231
rect 13860 29180 13877 29197
rect 7857 29146 7874 29163
rect 8938 29146 8955 29163
rect 10686 29146 10703 29163
rect 12342 29146 12359 29163
rect 14734 29146 14751 29163
rect 15700 29146 15717 29163
rect 6914 29044 6931 29061
rect 10364 29044 10381 29061
rect 11376 29044 11393 29061
rect 11882 29044 11899 29061
rect 13768 29044 13785 29061
rect 15148 29044 15165 29061
rect 16390 29044 16407 29061
rect 8823 29010 8840 29027
rect 15700 29010 15717 29027
rect 10410 28976 10427 28993
rect 11146 28976 11163 28993
rect 16298 28976 16315 28993
rect 4798 28942 4815 28959
rect 6730 28942 6747 28959
rect 6799 28942 6816 28959
rect 6868 28942 6885 28959
rect 6960 28942 6977 28959
rect 7420 28942 7437 28959
rect 7466 28942 7483 28959
rect 7512 28942 7529 28959
rect 8432 28942 8449 28959
rect 8524 28942 8541 28959
rect 8754 28942 8771 28959
rect 8892 28942 8909 28959
rect 8984 28942 9001 28959
rect 10272 28942 10289 28959
rect 10318 28942 10335 28959
rect 11192 28942 11209 28959
rect 11698 28942 11715 28959
rect 11790 28942 11807 28959
rect 13768 28942 13785 28959
rect 13860 28942 13877 28959
rect 14108 28942 14125 28959
rect 15148 28942 15165 28959
rect 15240 28942 15257 28959
rect 15792 28942 15809 28959
rect 15838 28942 15855 28959
rect 16206 28942 16223 28959
rect 16252 28942 16269 28959
rect 16390 28942 16407 28959
rect 17034 28942 17051 28959
rect 17080 28942 17097 28959
rect 17126 28942 17143 28959
rect 17448 28942 17465 28959
rect 17540 28942 17557 28959
rect 4936 28908 4953 28925
rect 8478 28908 8495 28925
rect 15700 28908 15717 28925
rect 17632 28908 17649 28925
rect 5672 28874 5689 28891
rect 8938 28874 8955 28891
rect 14159 28874 14176 28891
rect 17218 28874 17235 28891
rect 5580 28772 5597 28789
rect 6914 28772 6931 28789
rect 8846 28772 8863 28789
rect 15838 28772 15855 28789
rect 21036 28772 21053 28789
rect 6270 28738 6287 28755
rect 10318 28738 10335 28755
rect 18460 28738 18477 28755
rect 6592 28704 6609 28721
rect 6868 28704 6885 28721
rect 6960 28704 6977 28721
rect 7006 28704 7023 28721
rect 8110 28704 8127 28721
rect 8179 28704 8196 28721
rect 8340 28704 8357 28721
rect 8800 28704 8817 28721
rect 8892 28704 8909 28721
rect 10410 28704 10427 28721
rect 10456 28704 10473 28721
rect 13354 28704 13371 28721
rect 15792 28704 15809 28721
rect 15884 28704 15901 28721
rect 17126 28704 17143 28721
rect 4706 28670 4723 28687
rect 4844 28670 4861 28687
rect 6638 28670 6655 28687
rect 13400 28670 13417 28687
rect 13492 28670 13509 28687
rect 17080 28670 17097 28687
rect 17218 28670 17235 28687
rect 17448 28670 17465 28687
rect 17586 28670 17603 28687
rect 20162 28670 20179 28687
rect 20300 28670 20317 28687
rect 7006 28636 7023 28653
rect 8248 28636 8265 28653
rect 8294 28602 8311 28619
rect 10364 28602 10381 28619
rect 13446 28602 13463 28619
rect 17172 28602 17189 28619
rect 5166 28500 5183 28517
rect 20300 28500 20317 28517
rect 6868 28466 6885 28483
rect 16666 28466 16683 28483
rect 5488 28432 5505 28449
rect 12940 28432 12957 28449
rect 13952 28432 13969 28449
rect 15240 28432 15257 28449
rect 15700 28432 15717 28449
rect 15792 28432 15809 28449
rect 15930 28432 15947 28449
rect 15976 28432 15993 28449
rect 20576 28432 20593 28449
rect 5350 28398 5367 28415
rect 6684 28398 6701 28415
rect 6776 28398 6793 28415
rect 8432 28398 8449 28415
rect 10180 28398 10197 28415
rect 14228 28398 14245 28415
rect 16620 28398 16637 28415
rect 16728 28398 16745 28415
rect 17218 28398 17235 28415
rect 17346 28398 17363 28415
rect 19288 28398 19305 28415
rect 19702 28398 19719 28415
rect 20484 28398 20501 28415
rect 8592 28364 8609 28381
rect 8643 28364 8660 28381
rect 10303 28364 10320 28381
rect 13078 28364 13095 28381
rect 14366 28364 14383 28381
rect 19472 28364 19489 28381
rect 5396 28330 5413 28347
rect 9467 28330 9484 28347
rect 10870 28330 10887 28347
rect 16850 28330 16867 28347
rect 17908 28330 17925 28347
rect 19288 28330 19305 28347
rect 20530 28330 20547 28347
rect 5212 28228 5229 28245
rect 5396 28228 5413 28245
rect 8984 28228 9001 28245
rect 10548 28228 10565 28245
rect 10594 28228 10611 28245
rect 12894 28228 12911 28245
rect 14642 28228 14659 28245
rect 15470 28228 15487 28245
rect 17356 28228 17373 28245
rect 17770 28228 17787 28245
rect 19380 28228 19397 28245
rect 21082 28228 21099 28245
rect 9766 28194 9783 28211
rect 10226 28194 10243 28211
rect 11974 28194 11991 28211
rect 18138 28194 18155 28211
rect 5442 28160 5459 28177
rect 8800 28160 8817 28177
rect 8938 28160 8955 28177
rect 9030 28160 9047 28177
rect 9674 28160 9691 28177
rect 10134 28160 10151 28177
rect 10272 28160 10289 28177
rect 10510 28160 10527 28177
rect 11836 28160 11853 28177
rect 12020 28160 12037 28177
rect 12802 28160 12819 28177
rect 12894 28160 12911 28177
rect 13308 28160 13325 28177
rect 13400 28160 13417 28177
rect 14320 28160 14337 28177
rect 14367 28160 14384 28177
rect 14458 28160 14475 28177
rect 14504 28160 14521 28177
rect 14553 28160 14570 28177
rect 15470 28160 15487 28177
rect 15654 28160 15671 28177
rect 15838 28160 15855 28177
rect 17080 28160 17097 28177
rect 17218 28160 17235 28177
rect 17862 28160 17879 28177
rect 18092 28160 18109 28177
rect 18184 28160 18201 28177
rect 18824 28160 18841 28177
rect 5488 28126 5505 28143
rect 10686 28126 10703 28143
rect 11744 28126 11761 28143
rect 13354 28126 13371 28143
rect 17310 28126 17327 28143
rect 17816 28126 17833 28143
rect 18690 28126 18707 28143
rect 20208 28126 20225 28143
rect 20346 28126 20363 28143
rect 10134 28092 10151 28109
rect 17678 28092 17695 28109
rect 8869 28058 8886 28075
rect 10548 28058 10565 28075
rect 10456 27956 10473 27973
rect 17724 27956 17741 27973
rect 20346 27956 20363 27973
rect 17402 27922 17419 27939
rect 17172 27888 17189 27905
rect 17448 27888 17465 27905
rect 20622 27888 20639 27905
rect 10410 27854 10427 27871
rect 10502 27854 10519 27871
rect 11606 27854 11623 27871
rect 11698 27854 11715 27871
rect 12066 27854 12083 27871
rect 12388 27854 12405 27871
rect 17264 27854 17281 27871
rect 17678 27854 17695 27871
rect 17770 27854 17787 27871
rect 18690 27854 18707 27871
rect 19628 27854 19645 27871
rect 20530 27854 20547 27871
rect 17724 27820 17741 27837
rect 18813 27820 18830 27837
rect 11652 27786 11669 27803
rect 11974 27786 11991 27803
rect 19380 27786 19397 27803
rect 19679 27786 19696 27803
rect 20576 27786 20593 27803
rect 6776 27684 6793 27701
rect 4733 27650 4750 27667
rect 7374 27650 7391 27667
rect 11652 27650 11669 27667
rect 18414 27650 18431 27667
rect 18920 27650 18937 27667
rect 4683 27616 4700 27633
rect 6454 27616 6471 27633
rect 6546 27616 6563 27633
rect 6776 27616 6793 27633
rect 10272 27616 10289 27633
rect 10410 27616 10427 27633
rect 10456 27616 10473 27633
rect 11606 27616 11623 27633
rect 11698 27616 11715 27633
rect 11974 27616 11991 27633
rect 12112 27616 12129 27633
rect 12250 27616 12267 27633
rect 13354 27616 13371 27633
rect 13446 27616 13463 27633
rect 13492 27616 13509 27633
rect 15148 27616 15165 27633
rect 15286 27616 15303 27633
rect 15700 27616 15717 27633
rect 15792 27616 15809 27633
rect 18000 27616 18017 27633
rect 18092 27616 18109 27633
rect 18460 27616 18477 27633
rect 19012 27616 19029 27633
rect 4522 27582 4539 27599
rect 5557 27582 5574 27599
rect 6914 27582 6931 27599
rect 7328 27582 7345 27599
rect 12342 27582 12359 27599
rect 15378 27582 15395 27599
rect 15470 27582 15487 27599
rect 19104 27582 19121 27599
rect 6822 27548 6839 27565
rect 7190 27548 7207 27565
rect 15746 27548 15763 27565
rect 18322 27548 18339 27565
rect 6500 27514 6517 27531
rect 7236 27514 7253 27531
rect 13354 27514 13371 27531
rect 18046 27514 18063 27531
rect 18552 27514 18569 27531
rect 18736 27412 18753 27429
rect 20185 27412 20202 27429
rect 14964 27378 14981 27395
rect 6385 27344 6402 27361
rect 7558 27344 7575 27361
rect 7650 27344 7667 27361
rect 9536 27344 9553 27361
rect 18782 27344 18799 27361
rect 5350 27310 5367 27327
rect 5511 27310 5528 27327
rect 7512 27310 7529 27327
rect 7604 27310 7621 27327
rect 8662 27310 8679 27327
rect 8800 27310 8817 27327
rect 9352 27310 9369 27327
rect 9720 27310 9737 27327
rect 13124 27310 13141 27327
rect 13258 27310 13275 27327
rect 15102 27310 15119 27327
rect 16482 27310 16499 27327
rect 16574 27310 16591 27327
rect 18644 27310 18661 27327
rect 18690 27310 18707 27327
rect 19150 27310 19167 27327
rect 19311 27310 19328 27327
rect 5561 27276 5578 27293
rect 8754 27276 8771 27293
rect 14964 27276 14981 27293
rect 19361 27276 19378 27293
rect 7420 27242 7437 27259
rect 9306 27242 9323 27259
rect 13814 27242 13831 27259
rect 15056 27242 15073 27259
rect 16528 27242 16545 27259
rect 5557 27140 5574 27157
rect 6040 27140 6057 27157
rect 6270 27140 6287 27157
rect 7765 27140 7782 27157
rect 11928 27140 11945 27157
rect 13492 27140 13509 27157
rect 15286 27140 15303 27157
rect 18368 27140 18385 27157
rect 6937 27106 6954 27123
rect 8156 27106 8173 27123
rect 9398 27106 9415 27123
rect 10640 27106 10657 27123
rect 10740 27106 10757 27123
rect 14730 27106 14747 27123
rect 16390 27106 16407 27123
rect 4677 27072 4694 27089
rect 4721 27072 4738 27089
rect 6224 27072 6241 27089
rect 6730 27072 6747 27089
rect 6891 27072 6908 27089
rect 8248 27072 8265 27089
rect 8892 27072 8909 27089
rect 9260 27072 9277 27089
rect 11836 27072 11853 27089
rect 11974 27072 11991 27089
rect 12204 27072 12221 27089
rect 12296 27072 12313 27089
rect 16344 27072 16361 27089
rect 16482 27072 16499 27089
rect 4522 27038 4539 27055
rect 6270 27038 6287 27055
rect 6362 27038 6379 27055
rect 8938 27038 8955 27055
rect 8984 27038 9001 27055
rect 9398 27038 9415 27055
rect 13354 27038 13371 27055
rect 13400 27038 13417 27055
rect 13492 27038 13509 27055
rect 14596 27038 14613 27055
rect 16528 27038 16545 27055
rect 18230 27038 18247 27055
rect 18276 27038 18293 27055
rect 18368 27038 18385 27055
rect 20300 27038 20317 27055
rect 20438 27038 20455 27055
rect 21312 27038 21329 27055
rect 9306 27004 9323 27021
rect 11836 27004 11853 27021
rect 8340 26970 8357 26987
rect 8800 26970 8817 26987
rect 9352 26970 9369 26987
rect 10732 26970 10749 26987
rect 10824 26970 10841 26987
rect 12204 26970 12221 26987
rect 16574 26970 16591 26987
rect 17954 26868 17971 26885
rect 15056 26834 15073 26851
rect 6776 26800 6793 26817
rect 7604 26800 7621 26817
rect 7650 26800 7667 26817
rect 8662 26800 8679 26817
rect 16482 26800 16499 26817
rect 18000 26800 18017 26817
rect 6638 26766 6655 26783
rect 6960 26766 6977 26783
rect 7512 26766 7529 26783
rect 7558 26766 7575 26783
rect 10272 26766 10289 26783
rect 10406 26766 10423 26783
rect 11284 26766 11301 26783
rect 11418 26766 11435 26783
rect 12204 26766 12221 26783
rect 12296 26766 12313 26783
rect 14642 26766 14659 26783
rect 14872 26766 14889 26783
rect 14949 26766 14966 26783
rect 16616 26766 16633 26783
rect 17816 26766 17833 26783
rect 19150 26766 19167 26783
rect 7420 26732 7437 26749
rect 8524 26732 8541 26749
rect 19310 26732 19327 26749
rect 19361 26732 19378 26749
rect 8340 26698 8357 26715
rect 8570 26698 8587 26715
rect 10962 26698 10979 26715
rect 11974 26698 11991 26715
rect 12250 26698 12267 26715
rect 17172 26698 17189 26715
rect 17862 26698 17879 26715
rect 17908 26698 17925 26715
rect 20185 26698 20202 26715
rect 6270 26596 6287 26613
rect 6960 26596 6977 26613
rect 10732 26596 10749 26613
rect 20392 26596 20409 26613
rect 20622 26596 20639 26613
rect 11878 26562 11895 26579
rect 15792 26562 15809 26579
rect 15884 26562 15901 26579
rect 20576 26562 20593 26579
rect 21289 26562 21306 26579
rect 6224 26528 6241 26545
rect 6960 26528 6977 26545
rect 7052 26528 7069 26545
rect 7190 26528 7207 26545
rect 7282 26528 7299 26545
rect 9260 26528 9277 26545
rect 10548 26528 10565 26545
rect 11744 26528 11761 26545
rect 13492 26528 13509 26545
rect 13538 26528 13555 26545
rect 13676 26528 13693 26545
rect 15194 26528 15211 26545
rect 15930 26528 15947 26545
rect 16252 26528 16269 26545
rect 17816 26528 17833 26545
rect 18230 26528 18247 26545
rect 18322 26528 18339 26545
rect 21243 26528 21260 26545
rect 6270 26494 6287 26511
rect 6362 26494 6379 26511
rect 9306 26494 9323 26511
rect 9352 26494 9369 26511
rect 10502 26494 10519 26511
rect 13584 26494 13601 26511
rect 15148 26494 15165 26511
rect 15378 26494 15395 26511
rect 16206 26494 16223 26511
rect 17770 26494 17787 26511
rect 18000 26494 18017 26511
rect 20668 26494 20685 26511
rect 21082 26494 21099 26511
rect 18230 26460 18247 26477
rect 6040 26426 6057 26443
rect 9076 26426 9093 26443
rect 12434 26426 12451 26443
rect 13676 26426 13693 26443
rect 15930 26426 15947 26443
rect 16390 26426 16407 26443
rect 22117 26426 22134 26443
rect 6569 26324 6586 26341
rect 12112 26324 12129 26341
rect 16344 26324 16361 26341
rect 17862 26324 17879 26341
rect 8018 26256 8035 26273
rect 8110 26256 8127 26273
rect 13308 26256 13325 26273
rect 13630 26256 13647 26273
rect 14964 26256 14981 26273
rect 5534 26222 5551 26239
rect 5695 26222 5712 26239
rect 8432 26222 8449 26239
rect 8587 26222 8604 26239
rect 11606 26222 11623 26239
rect 11698 26222 11715 26239
rect 12112 26222 12129 26239
rect 12204 26222 12221 26239
rect 12940 26222 12957 26239
rect 13262 26222 13279 26239
rect 13758 26222 13775 26239
rect 14780 26222 14797 26239
rect 15056 26222 15073 26239
rect 16298 26222 16315 26239
rect 16344 26222 16361 26239
rect 17908 26222 17925 26239
rect 19104 26222 19121 26239
rect 5741 26188 5758 26205
rect 7972 26188 7989 26205
rect 8631 26188 8648 26205
rect 11652 26188 11669 26205
rect 16206 26188 16223 26205
rect 17724 26188 17741 26205
rect 17954 26188 17971 26205
rect 19264 26188 19281 26205
rect 19311 26188 19328 26205
rect 20139 26188 20156 26205
rect 6569 26154 6586 26171
rect 7788 26154 7805 26171
rect 9467 26154 9484 26171
rect 14320 26154 14337 26171
rect 16436 26154 16453 26171
rect 17770 26154 17787 26171
rect 6914 26052 6931 26069
rect 13768 26052 13785 26069
rect 18506 26052 18523 26069
rect 4637 26018 4654 26035
rect 7493 26018 7510 26035
rect 9236 26018 9253 26035
rect 17950 26018 17967 26035
rect 20415 26018 20432 26035
rect 21496 26018 21513 26035
rect 23244 26018 23261 26035
rect 4591 25984 4608 26001
rect 6868 25984 6885 26001
rect 7443 25984 7460 26001
rect 9275 25984 9292 26001
rect 12940 25984 12957 26001
rect 13262 25984 13279 26001
rect 13400 25984 13417 26001
rect 13630 25984 13647 26001
rect 17816 25984 17833 26001
rect 20369 25984 20386 26001
rect 21680 25984 21697 26001
rect 23106 25984 23123 26001
rect 23152 25984 23169 26001
rect 23290 25984 23307 26001
rect 23336 25984 23353 26001
rect 4430 25950 4447 25967
rect 7006 25950 7023 25967
rect 7282 25950 7299 25967
rect 9076 25950 9093 25967
rect 13676 25950 13693 25967
rect 13768 25950 13785 25967
rect 20208 25950 20225 25967
rect 21531 25950 21548 25967
rect 21588 25950 21605 25967
rect 23382 25950 23399 25967
rect 5465 25882 5482 25899
rect 6684 25882 6701 25899
rect 8317 25882 8334 25899
rect 10111 25882 10128 25899
rect 13078 25882 13095 25899
rect 21243 25882 21260 25899
rect 21634 25882 21651 25899
rect 9076 25780 9093 25797
rect 16390 25780 16407 25797
rect 17494 25780 17511 25797
rect 23014 25780 23031 25797
rect 8984 25746 9001 25763
rect 9168 25712 9185 25729
rect 13722 25712 13739 25729
rect 16160 25712 16177 25729
rect 17264 25712 17281 25729
rect 23060 25712 23077 25729
rect 4660 25678 4677 25695
rect 4815 25678 4832 25695
rect 4859 25678 4876 25695
rect 7742 25678 7759 25695
rect 7834 25678 7851 25695
rect 8248 25678 8265 25695
rect 8340 25678 8357 25695
rect 8524 25678 8541 25695
rect 8754 25678 8771 25695
rect 9122 25678 9139 25695
rect 13676 25678 13693 25695
rect 13768 25678 13785 25695
rect 16206 25678 16223 25695
rect 17310 25678 17327 25695
rect 20576 25678 20593 25695
rect 21588 25678 21605 25695
rect 22830 25678 22847 25695
rect 22876 25678 22893 25695
rect 23106 25678 23123 25695
rect 7788 25644 7805 25661
rect 8984 25644 9001 25661
rect 5695 25610 5712 25627
rect 20622 25610 20639 25627
rect 21634 25610 21651 25627
rect 7535 25508 7552 25525
rect 8064 25508 8081 25525
rect 18874 25508 18891 25525
rect 23658 25508 23675 25525
rect 6711 25474 6728 25491
rect 19196 25474 19213 25491
rect 3372 25440 3389 25457
rect 3527 25440 3544 25457
rect 3571 25440 3588 25457
rect 6500 25440 6517 25457
rect 6655 25440 6672 25457
rect 8064 25440 8081 25457
rect 9829 25440 9846 25457
rect 9873 25440 9890 25457
rect 18690 25440 18707 25457
rect 19104 25440 19121 25457
rect 19242 25440 19259 25457
rect 23520 25440 23537 25457
rect 8202 25406 8219 25423
rect 9674 25406 9691 25423
rect 18736 25406 18753 25423
rect 23428 25406 23445 25423
rect 23704 25406 23721 25423
rect 8110 25372 8127 25389
rect 4407 25338 4424 25355
rect 10709 25338 10726 25355
rect 19104 25338 19121 25355
rect 23566 25338 23583 25355
rect 17402 25236 17419 25253
rect 22715 25236 22732 25253
rect 3142 25168 3159 25185
rect 17172 25168 17189 25185
rect 18506 25168 18523 25185
rect 20392 25168 20409 25185
rect 3297 25134 3314 25151
rect 4177 25134 4194 25151
rect 4660 25134 4677 25151
rect 4798 25134 4815 25151
rect 4844 25134 4861 25151
rect 8662 25134 8679 25151
rect 11008 25134 11025 25151
rect 11169 25134 11186 25151
rect 14872 25134 14889 25151
rect 14918 25134 14935 25151
rect 14964 25134 14981 25151
rect 17218 25134 17235 25151
rect 17770 25134 17787 25151
rect 18640 25134 18657 25151
rect 20346 25134 20363 25151
rect 21680 25134 21697 25151
rect 21841 25134 21858 25151
rect 3353 25100 3370 25117
rect 4752 25100 4769 25117
rect 8822 25100 8839 25117
rect 8873 25100 8890 25117
rect 11219 25100 11236 25117
rect 17632 25100 17649 25117
rect 17724 25100 17741 25117
rect 21891 25100 21908 25117
rect 4936 25066 4953 25083
rect 9697 25066 9714 25083
rect 12043 25066 12060 25083
rect 15056 25066 15073 25083
rect 17770 25066 17787 25083
rect 19196 25066 19213 25083
rect 20530 25066 20547 25083
rect 12894 24964 12911 24981
rect 9827 24930 9844 24947
rect 11771 24930 11788 24947
rect 6040 24896 6057 24913
rect 6097 24896 6114 24913
rect 6191 24896 6208 24913
rect 6246 24891 6263 24908
rect 6301 24896 6318 24913
rect 6352 24896 6369 24913
rect 9783 24896 9800 24913
rect 11715 24896 11732 24913
rect 12986 24896 13003 24913
rect 13124 24896 13141 24913
rect 13262 24896 13279 24913
rect 13354 24896 13371 24913
rect 14872 24896 14889 24913
rect 15148 24896 15165 24913
rect 15194 24896 15211 24913
rect 15332 24896 15349 24913
rect 15838 24896 15855 24913
rect 15884 24896 15901 24913
rect 15930 24896 15947 24913
rect 17080 24896 17097 24913
rect 17356 24896 17373 24913
rect 18276 24896 18293 24913
rect 18736 24896 18753 24913
rect 20346 24896 20363 24913
rect 21404 24896 21421 24913
rect 9628 24862 9645 24879
rect 11560 24862 11577 24879
rect 18322 24862 18339 24879
rect 18414 24862 18431 24879
rect 18690 24862 18707 24879
rect 18920 24862 18937 24879
rect 20392 24862 20409 24879
rect 21450 24862 21467 24879
rect 18368 24828 18385 24845
rect 21588 24828 21605 24845
rect 6040 24794 6057 24811
rect 10663 24794 10680 24811
rect 12595 24794 12612 24811
rect 13400 24794 13417 24811
rect 14872 24794 14889 24811
rect 16022 24794 16039 24811
rect 17126 24794 17143 24811
rect 20484 24794 20501 24811
rect 6569 24692 6586 24709
rect 18690 24692 18707 24709
rect 22991 24692 23008 24709
rect 24026 24692 24043 24709
rect 15838 24658 15855 24675
rect 7742 24624 7759 24641
rect 14780 24624 14797 24641
rect 15010 24624 15027 24641
rect 15056 24624 15073 24641
rect 18598 24624 18615 24641
rect 5534 24590 5551 24607
rect 5689 24590 5706 24607
rect 7929 24590 7946 24607
rect 8202 24590 8219 24607
rect 8401 24590 8418 24607
rect 10502 24590 10519 24607
rect 10559 24590 10576 24607
rect 10653 24588 10670 24605
rect 10709 24596 10726 24613
rect 10763 24596 10780 24613
rect 10814 24590 10831 24607
rect 11100 24590 11117 24607
rect 11261 24590 11278 24607
rect 13032 24590 13049 24607
rect 13308 24590 13325 24607
rect 13768 24590 13785 24607
rect 13952 24590 13969 24607
rect 14044 24590 14061 24607
rect 16712 24590 16729 24607
rect 16942 24590 16959 24607
rect 17080 24590 17097 24607
rect 17218 24590 17235 24607
rect 18552 24590 18569 24607
rect 19564 24590 19581 24607
rect 19763 24590 19780 24607
rect 21956 24590 21973 24607
rect 23980 24590 23997 24607
rect 5745 24556 5762 24573
rect 7742 24556 7759 24573
rect 7834 24556 7851 24573
rect 7880 24556 7897 24573
rect 8362 24556 8379 24573
rect 11311 24556 11328 24573
rect 15746 24556 15763 24573
rect 19724 24556 19741 24573
rect 22116 24556 22133 24573
rect 22167 24556 22184 24573
rect 24072 24556 24089 24573
rect 9237 24522 9254 24539
rect 10732 24522 10749 24539
rect 12135 24522 12152 24539
rect 13078 24522 13095 24539
rect 13676 24522 13693 24539
rect 14872 24522 14889 24539
rect 16620 24522 16637 24539
rect 20599 24522 20616 24539
rect 7949 24420 7966 24437
rect 17770 24420 17787 24437
rect 23428 24420 23445 24437
rect 9306 24386 9323 24403
rect 23484 24386 23501 24403
rect 24302 24386 24319 24403
rect 3619 24352 3636 24369
rect 3663 24352 3680 24369
rect 7069 24352 7086 24369
rect 7113 24352 7130 24369
rect 9168 24352 9185 24369
rect 9260 24352 9277 24369
rect 9355 24352 9372 24369
rect 12020 24352 12037 24369
rect 12077 24352 12094 24369
rect 12171 24352 12188 24369
rect 12233 24347 12250 24364
rect 12281 24347 12298 24364
rect 12332 24352 12349 24369
rect 16068 24352 16085 24369
rect 16160 24352 16177 24369
rect 16344 24352 16361 24369
rect 17586 24352 17603 24369
rect 20346 24352 20363 24369
rect 20760 24352 20777 24369
rect 20898 24352 20915 24369
rect 20990 24352 21007 24369
rect 21128 24352 21145 24369
rect 22968 24352 22985 24369
rect 23382 24352 23399 24369
rect 23934 24352 23951 24369
rect 24026 24352 24043 24369
rect 24072 24352 24089 24369
rect 3464 24318 3481 24335
rect 6914 24318 6931 24335
rect 9306 24318 9323 24335
rect 17540 24318 17557 24335
rect 20392 24318 20409 24335
rect 20530 24318 20547 24335
rect 21174 24318 21191 24335
rect 22922 24318 22939 24335
rect 23566 24318 23583 24335
rect 16344 24284 16361 24301
rect 23152 24284 23169 24301
rect 24348 24284 24365 24301
rect 4499 24250 4516 24267
rect 12020 24250 12037 24267
rect 23428 24250 23445 24267
rect 23934 24250 23951 24267
rect 9099 24148 9116 24165
rect 22761 24148 22778 24165
rect 5028 24114 5045 24131
rect 18460 24114 18477 24131
rect 20668 24114 20685 24131
rect 24486 24114 24503 24131
rect 3142 24080 3159 24097
rect 8064 24080 8081 24097
rect 12342 24080 12359 24097
rect 17080 24080 17097 24097
rect 20438 24080 20455 24097
rect 21726 24080 21743 24097
rect 24256 24080 24273 24097
rect 3303 24046 3320 24063
rect 5120 24046 5137 24063
rect 8225 24046 8242 24063
rect 12158 24046 12175 24063
rect 12296 24046 12313 24063
rect 12388 24046 12405 24063
rect 13998 24046 14015 24063
rect 14182 24046 14199 24063
rect 14274 24046 14291 24063
rect 16344 24046 16361 24063
rect 16850 24046 16867 24063
rect 17034 24046 17051 24063
rect 18598 24046 18615 24063
rect 20484 24046 20501 24063
rect 21887 24046 21904 24063
rect 24118 24046 24135 24063
rect 24164 24046 24181 24063
rect 24624 24046 24641 24063
rect 3353 24012 3370 24029
rect 4982 24012 4999 24029
rect 5074 24012 5091 24029
rect 8271 24012 8288 24029
rect 18460 24012 18477 24029
rect 21937 24012 21954 24029
rect 24256 24012 24273 24029
rect 24486 24012 24503 24029
rect 4177 23978 4194 23995
rect 13906 23978 13923 23995
rect 16390 23978 16407 23995
rect 16988 23978 17005 23995
rect 18552 23978 18569 23995
rect 24578 23978 24595 23995
rect 4982 23876 4999 23893
rect 19012 23876 19029 23893
rect 21404 23876 21421 23893
rect 23750 23876 23767 23893
rect 3624 23842 3641 23859
rect 3675 23842 3692 23859
rect 6362 23842 6379 23859
rect 7113 23842 7130 23859
rect 18456 23842 18473 23859
rect 21312 23842 21329 23859
rect 24103 23842 24120 23859
rect 4752 23808 4769 23825
rect 4819 23808 4836 23825
rect 4910 23808 4927 23825
rect 4965 23803 4982 23820
rect 5013 23808 5030 23825
rect 5064 23808 5081 23825
rect 6454 23808 6471 23825
rect 6500 23808 6517 23825
rect 6914 23808 6931 23825
rect 7074 23808 7091 23825
rect 9030 23808 9047 23825
rect 9185 23808 9202 23825
rect 9229 23808 9246 23825
rect 12986 23808 13003 23825
rect 13078 23808 13095 23825
rect 14964 23808 14981 23825
rect 15056 23808 15073 23825
rect 17908 23808 17925 23825
rect 18322 23808 18339 23825
rect 21450 23808 21467 23825
rect 23980 23808 23997 23825
rect 3464 23774 3481 23791
rect 4499 23774 4516 23791
rect 7949 23774 7966 23791
rect 13216 23774 13233 23791
rect 15194 23774 15211 23791
rect 17954 23774 17971 23791
rect 18092 23774 18109 23791
rect 23612 23774 23629 23791
rect 23658 23774 23675 23791
rect 23750 23774 23767 23791
rect 6362 23706 6379 23723
rect 10065 23706 10082 23723
rect 21312 23706 21329 23723
rect 24670 23706 24687 23723
rect 6684 23604 6701 23621
rect 18552 23604 18569 23621
rect 20415 23604 20432 23621
rect 6408 23570 6425 23587
rect 21220 23570 21237 23587
rect 9490 23536 9507 23553
rect 17862 23536 17879 23553
rect 18460 23536 18477 23553
rect 18598 23536 18615 23553
rect 19380 23536 19397 23553
rect 21818 23536 21835 23553
rect 22853 23536 22870 23553
rect 23152 23536 23169 23553
rect 5120 23502 5137 23519
rect 5281 23502 5298 23519
rect 6546 23502 6563 23519
rect 8156 23502 8173 23519
rect 8311 23502 8328 23519
rect 9444 23502 9461 23519
rect 9536 23502 9553 23519
rect 10180 23502 10197 23519
rect 10226 23502 10243 23519
rect 10318 23502 10335 23519
rect 10410 23502 10427 23519
rect 11008 23502 11025 23519
rect 11207 23502 11224 23519
rect 12986 23502 13003 23519
rect 13262 23502 13279 23519
rect 17678 23502 17695 23519
rect 17770 23502 17787 23519
rect 17908 23502 17925 23519
rect 18506 23502 18523 23519
rect 19541 23502 19558 23519
rect 21358 23502 21375 23519
rect 21979 23502 21996 23519
rect 23198 23502 23215 23519
rect 24302 23502 24319 23519
rect 24436 23502 24453 23519
rect 5331 23468 5348 23485
rect 8367 23468 8384 23485
rect 10364 23468 10381 23485
rect 11168 23468 11185 23485
rect 19587 23468 19604 23485
rect 21220 23468 21237 23485
rect 22029 23468 22046 23485
rect 6155 23434 6172 23451
rect 6500 23434 6517 23451
rect 6592 23434 6609 23451
rect 9191 23434 9208 23451
rect 10272 23434 10289 23451
rect 12043 23434 12060 23451
rect 13032 23434 13049 23451
rect 21312 23434 21329 23451
rect 23382 23434 23399 23451
rect 24992 23434 25009 23451
rect 10249 23332 10266 23349
rect 10686 23332 10703 23349
rect 10732 23332 10749 23349
rect 10824 23332 10841 23349
rect 14642 23332 14659 23349
rect 17126 23332 17143 23349
rect 17954 23332 17971 23349
rect 6270 23298 6287 23315
rect 6362 23298 6379 23315
rect 9421 23298 9438 23315
rect 12020 23298 12037 23315
rect 12112 23298 12129 23315
rect 20572 23298 20589 23315
rect 21492 23298 21509 23315
rect 6408 23264 6425 23281
rect 6472 23264 6489 23281
rect 9369 23264 9386 23281
rect 10640 23264 10657 23281
rect 11560 23264 11577 23281
rect 11652 23264 11669 23281
rect 12158 23264 12175 23281
rect 12214 23264 12231 23281
rect 13124 23264 13141 23281
rect 13262 23264 13279 23281
rect 14734 23264 14751 23281
rect 14872 23264 14889 23281
rect 16298 23264 16315 23281
rect 16528 23264 16545 23281
rect 17126 23264 17143 23281
rect 17218 23264 17235 23281
rect 17908 23264 17925 23281
rect 18138 23264 18155 23281
rect 19012 23264 19029 23281
rect 19288 23264 19305 23281
rect 19380 23264 19397 23281
rect 21358 23264 21375 23281
rect 6316 23230 6333 23247
rect 9214 23230 9231 23247
rect 10824 23230 10841 23247
rect 11606 23230 11623 23247
rect 12066 23230 12083 23247
rect 13216 23230 13233 23247
rect 14964 23230 14981 23247
rect 16574 23230 16591 23247
rect 17310 23230 17327 23247
rect 20438 23230 20455 23247
rect 21128 23162 21145 23179
rect 22048 23162 22065 23179
rect 6523 23060 6540 23077
rect 9352 23060 9369 23077
rect 12135 23060 12152 23077
rect 16666 23060 16683 23077
rect 17540 23060 17557 23077
rect 21312 23060 21329 23077
rect 21680 23060 21697 23077
rect 22692 23060 22709 23077
rect 19886 23026 19903 23043
rect 15102 22992 15119 23009
rect 17862 22992 17879 23009
rect 17954 22992 17971 23009
rect 19656 22992 19673 23009
rect 20208 22992 20225 23009
rect 21220 22992 21237 23009
rect 21358 22992 21375 23009
rect 21726 22992 21743 23009
rect 5488 22958 5505 22975
rect 9306 22958 9323 22975
rect 9398 22958 9415 22975
rect 11100 22958 11117 22975
rect 11261 22958 11278 22975
rect 13354 22958 13371 22975
rect 13630 22958 13647 22975
rect 14964 22958 14981 22975
rect 15056 22958 15073 22975
rect 16114 22958 16131 22975
rect 16252 22958 16269 22975
rect 16666 22958 16683 22975
rect 16896 22958 16913 22975
rect 17494 22958 17511 22975
rect 17586 22958 17603 22975
rect 17816 22958 17833 22975
rect 19702 22958 19719 22975
rect 20346 22958 20363 22975
rect 21266 22958 21283 22975
rect 21588 22958 21605 22975
rect 21634 22958 21651 22975
rect 22462 22958 22479 22975
rect 22968 22958 22985 22975
rect 23060 22958 23077 22975
rect 24624 22958 24641 22975
rect 5648 22924 5665 22941
rect 5699 22924 5716 22941
rect 11307 22924 11324 22941
rect 13722 22924 13739 22941
rect 22738 22924 22755 22941
rect 24784 22924 24801 22941
rect 24835 22924 24852 22941
rect 13400 22890 13417 22907
rect 16114 22890 16131 22907
rect 17954 22890 17971 22907
rect 20668 22890 20685 22907
rect 23014 22890 23031 22907
rect 25659 22890 25676 22907
rect 11077 22788 11094 22805
rect 14688 22788 14705 22805
rect 18322 22788 18339 22805
rect 19380 22788 19397 22805
rect 28419 22754 28436 22771
rect 3573 22720 3590 22737
rect 3617 22720 3634 22737
rect 7437 22720 7454 22737
rect 7481 22720 7498 22737
rect 10197 22720 10214 22737
rect 10241 22720 10258 22737
rect 12940 22720 12957 22737
rect 13032 22720 13049 22737
rect 13400 22720 13417 22737
rect 13630 22720 13647 22737
rect 14780 22720 14797 22737
rect 14872 22720 14889 22737
rect 15746 22720 15763 22737
rect 15884 22720 15901 22737
rect 15976 22720 15993 22737
rect 17766 22720 17783 22737
rect 19196 22720 19213 22737
rect 20070 22720 20087 22737
rect 23372 22720 23389 22737
rect 24210 22720 24227 22737
rect 28367 22720 28384 22737
rect 3418 22686 3435 22703
rect 7282 22686 7299 22703
rect 10042 22686 10059 22703
rect 13078 22686 13095 22703
rect 13676 22686 13693 22703
rect 16022 22686 16039 22703
rect 17632 22686 17649 22703
rect 18552 22686 18569 22703
rect 18598 22686 18615 22703
rect 18690 22686 18707 22703
rect 19242 22686 19259 22703
rect 20116 22686 20133 22703
rect 23244 22686 23261 22703
rect 24164 22686 24181 22703
rect 24302 22686 24319 22703
rect 28212 22686 28229 22703
rect 20254 22652 20271 22669
rect 23934 22652 23951 22669
rect 4453 22618 4470 22635
rect 8317 22618 8334 22635
rect 18644 22618 18661 22635
rect 24256 22618 24273 22635
rect 29247 22618 29264 22635
rect 6339 22516 6356 22533
rect 8708 22516 8725 22533
rect 17816 22516 17833 22533
rect 19150 22516 19167 22533
rect 23290 22516 23307 22533
rect 8455 22448 8472 22465
rect 17724 22448 17741 22465
rect 18460 22448 18477 22465
rect 24394 22448 24411 22465
rect 3142 22414 3159 22431
rect 3297 22414 3314 22431
rect 4177 22414 4194 22431
rect 4660 22414 4677 22431
rect 4737 22414 4754 22431
rect 4811 22414 4828 22431
rect 4873 22404 4890 22421
rect 4921 22404 4938 22421
rect 4972 22414 4989 22431
rect 5304 22414 5321 22431
rect 5465 22414 5482 22431
rect 7420 22414 7437 22431
rect 7575 22414 7592 22431
rect 8708 22414 8725 22431
rect 8765 22414 8782 22431
rect 8859 22414 8876 22431
rect 8921 22404 8938 22421
rect 8969 22414 8986 22431
rect 9020 22414 9037 22431
rect 13400 22414 13417 22431
rect 13676 22414 13693 22431
rect 14780 22414 14797 22431
rect 14918 22414 14935 22431
rect 15056 22414 15073 22431
rect 16298 22414 16315 22431
rect 16436 22414 16453 22431
rect 17632 22414 17649 22431
rect 17816 22414 17833 22431
rect 21312 22414 21329 22431
rect 21473 22414 21490 22431
rect 22968 22414 22985 22431
rect 23060 22414 23077 22431
rect 23290 22414 23307 22431
rect 23382 22414 23399 22431
rect 24549 22414 24566 22431
rect 3341 22380 3358 22397
rect 5515 22380 5532 22397
rect 7631 22380 7648 22397
rect 18583 22380 18600 22397
rect 21523 22380 21540 22397
rect 24601 22380 24618 22397
rect 4660 22346 4677 22363
rect 13446 22346 13463 22363
rect 14826 22346 14843 22363
rect 16206 22346 16223 22363
rect 17678 22346 17695 22363
rect 22347 22346 22364 22363
rect 23014 22346 23031 22363
rect 25429 22346 25446 22363
rect 4545 22244 4562 22261
rect 8271 22244 8288 22261
rect 14964 22244 14981 22261
rect 16206 22244 16223 22261
rect 23980 22244 23997 22261
rect 7443 22210 7460 22227
rect 9329 22210 9346 22227
rect 18506 22210 18523 22227
rect 21293 22210 21310 22227
rect 23413 22210 23430 22227
rect 24348 22210 24365 22227
rect 25544 22210 25561 22227
rect 26395 22210 26412 22227
rect 28469 22210 28486 22227
rect 3665 22176 3682 22193
rect 3709 22176 3726 22193
rect 7391 22176 7408 22193
rect 9122 22176 9139 22193
rect 9283 22176 9300 22193
rect 14964 22176 14981 22193
rect 15148 22176 15165 22193
rect 16206 22176 16223 22193
rect 16344 22176 16361 22193
rect 17632 22176 17649 22193
rect 17954 22176 17971 22193
rect 18092 22176 18109 22193
rect 18598 22176 18615 22193
rect 18644 22176 18661 22193
rect 21082 22176 21099 22193
rect 21243 22176 21260 22193
rect 23290 22176 23307 22193
rect 24256 22176 24273 22193
rect 25406 22176 25423 22193
rect 25498 22176 25515 22193
rect 25590 22176 25607 22193
rect 26349 22176 26366 22193
rect 28258 22176 28275 22193
rect 28413 22176 28430 22193
rect 3510 22142 3527 22159
rect 7236 22142 7253 22159
rect 16390 22142 16407 22159
rect 17770 22142 17787 22159
rect 24210 22142 24227 22159
rect 24348 22142 24365 22159
rect 26188 22142 26205 22159
rect 18506 22108 18523 22125
rect 10157 22074 10174 22091
rect 22117 22074 22134 22091
rect 25682 22074 25699 22091
rect 27223 22074 27240 22091
rect 29293 22074 29310 22091
rect 17678 21972 17695 21989
rect 23244 21972 23261 21989
rect 28028 21972 28045 21989
rect 25728 21938 25745 21955
rect 27775 21938 27792 21955
rect 6201 21904 6218 21921
rect 17080 21904 17097 21921
rect 17908 21904 17925 21921
rect 19518 21904 19535 21921
rect 21220 21904 21237 21921
rect 22255 21904 22272 21921
rect 24440 21904 24457 21921
rect 5166 21870 5183 21887
rect 5327 21870 5344 21887
rect 6454 21870 6471 21887
rect 6500 21870 6517 21887
rect 6592 21870 6609 21887
rect 6684 21870 6701 21887
rect 10180 21870 10197 21887
rect 10272 21870 10289 21887
rect 10318 21870 10335 21887
rect 10364 21870 10381 21887
rect 11330 21870 11347 21887
rect 11485 21870 11502 21887
rect 14412 21870 14429 21887
rect 14550 21870 14567 21887
rect 14964 21870 14981 21887
rect 15148 21870 15165 21887
rect 16344 21870 16361 21887
rect 16482 21870 16499 21887
rect 16528 21870 16545 21887
rect 16896 21870 16913 21887
rect 17034 21870 17051 21887
rect 17540 21870 17557 21887
rect 17862 21870 17879 21887
rect 19679 21870 19696 21887
rect 21381 21870 21398 21887
rect 22508 21870 22525 21887
rect 22565 21870 22582 21887
rect 22659 21870 22676 21887
rect 22707 21860 22724 21877
rect 22755 21860 22772 21877
rect 22820 21870 22837 21887
rect 23244 21870 23261 21887
rect 23336 21870 23353 21887
rect 25728 21870 25745 21887
rect 25866 21870 25883 21887
rect 26740 21870 26757 21887
rect 26895 21870 26912 21887
rect 28028 21870 28045 21887
rect 28085 21870 28102 21887
rect 28186 21870 28203 21887
rect 28234 21860 28251 21877
rect 28281 21876 28298 21893
rect 28340 21870 28357 21887
rect 5373 21836 5390 21853
rect 6638 21836 6655 21853
rect 11541 21836 11558 21853
rect 19729 21836 19746 21853
rect 21431 21836 21448 21853
rect 24600 21836 24617 21853
rect 24651 21836 24668 21853
rect 26951 21836 26968 21853
rect 6546 21802 6563 21819
rect 10456 21802 10473 21819
rect 12365 21802 12382 21819
rect 14320 21802 14337 21819
rect 14918 21802 14935 21819
rect 16344 21802 16361 21819
rect 16896 21802 16913 21819
rect 20553 21802 20570 21819
rect 22508 21802 22525 21819
rect 25475 21802 25492 21819
rect 25820 21802 25837 21819
rect 4798 21700 4815 21717
rect 18230 21700 18247 21717
rect 27177 21700 27194 21717
rect 3629 21666 3646 21683
rect 4752 21666 4769 21683
rect 7442 21666 7459 21683
rect 7493 21666 7510 21683
rect 9885 21666 9902 21683
rect 11863 21666 11880 21683
rect 13308 21666 13325 21683
rect 14531 21666 14548 21683
rect 17724 21666 17741 21683
rect 26353 21666 26370 21683
rect 28423 21666 28440 21683
rect 29247 21666 29264 21683
rect 3573 21632 3590 21649
rect 4844 21632 4861 21649
rect 4890 21632 4907 21649
rect 6408 21632 6425 21649
rect 6500 21632 6517 21649
rect 6638 21632 6655 21649
rect 9674 21632 9691 21649
rect 9829 21632 9846 21649
rect 11807 21632 11824 21649
rect 13032 21632 13049 21649
rect 13078 21632 13095 21649
rect 14475 21632 14492 21649
rect 15838 21632 15855 21649
rect 15884 21632 15901 21649
rect 16022 21632 16039 21649
rect 16160 21632 16177 21649
rect 16252 21632 16269 21649
rect 17494 21632 17511 21649
rect 17816 21632 17833 21649
rect 17954 21632 17971 21649
rect 18184 21632 18201 21649
rect 18322 21632 18339 21649
rect 26303 21632 26320 21649
rect 28212 21632 28229 21649
rect 28367 21632 28384 21649
rect 29500 21632 29517 21649
rect 29557 21632 29574 21649
rect 29658 21632 29675 21649
rect 29713 21627 29730 21644
rect 29761 21627 29778 21644
rect 29812 21632 29829 21649
rect 3418 21598 3435 21615
rect 7282 21598 7299 21615
rect 11652 21598 11669 21615
rect 14320 21598 14337 21615
rect 15355 21598 15372 21615
rect 18414 21598 18431 21615
rect 26142 21598 26159 21615
rect 12940 21564 12957 21581
rect 15654 21564 15671 21581
rect 4453 21530 4470 21547
rect 6454 21530 6471 21547
rect 8317 21530 8334 21547
rect 10709 21530 10726 21547
rect 12687 21530 12704 21547
rect 29500 21530 29517 21547
rect 6339 21428 6356 21445
rect 8110 21428 8127 21445
rect 9697 21428 9714 21445
rect 16620 21428 16637 21445
rect 20369 21394 20386 21411
rect 4798 21360 4815 21377
rect 10870 21360 10887 21377
rect 15217 21360 15234 21377
rect 19334 21360 19351 21377
rect 4862 21326 4879 21343
rect 5304 21326 5321 21343
rect 5465 21326 5482 21343
rect 8110 21326 8127 21343
rect 8187 21326 8204 21343
rect 8271 21326 8288 21343
rect 8317 21326 8334 21343
rect 8371 21316 8388 21333
rect 8422 21326 8439 21343
rect 8662 21326 8679 21343
rect 10594 21326 10611 21343
rect 10640 21326 10657 21343
rect 10778 21326 10795 21343
rect 10824 21326 10841 21343
rect 11422 21326 11439 21343
rect 14182 21326 14199 21343
rect 16390 21326 16407 21343
rect 16850 21326 16867 21343
rect 19495 21326 19512 21343
rect 4660 21292 4677 21309
rect 4752 21292 4769 21309
rect 4798 21292 4815 21309
rect 5515 21292 5532 21309
rect 8822 21292 8839 21309
rect 8873 21292 8890 21309
rect 10732 21292 10749 21309
rect 11582 21292 11599 21309
rect 11633 21292 11650 21309
rect 14342 21292 14359 21309
rect 14393 21292 14410 21309
rect 19545 21292 19562 21309
rect 12457 21258 12474 21275
rect 6500 21156 6517 21173
rect 8317 21156 8334 21173
rect 10571 21156 10588 21173
rect 12388 21156 12405 21173
rect 3721 21122 3738 21139
rect 6638 21122 6655 21139
rect 7442 21122 7459 21139
rect 7493 21122 7510 21139
rect 9747 21122 9764 21139
rect 18533 21122 18550 21139
rect 19357 21122 19374 21139
rect 23635 21122 23652 21139
rect 26027 21122 26044 21139
rect 3510 21088 3527 21105
rect 3671 21088 3688 21105
rect 4545 21088 4562 21105
rect 4798 21088 4815 21105
rect 4890 21088 4907 21105
rect 4936 21088 4953 21105
rect 5000 21088 5017 21105
rect 6500 21088 6517 21105
rect 6546 21088 6563 21105
rect 6684 21088 6701 21105
rect 6730 21088 6747 21105
rect 9697 21088 9714 21105
rect 12388 21088 12405 21105
rect 12445 21088 12462 21105
rect 12546 21088 12563 21105
rect 12601 21099 12618 21116
rect 12649 21099 12666 21116
rect 12700 21088 12717 21105
rect 18483 21088 18500 21105
rect 20116 21088 20133 21105
rect 20173 21088 20190 21105
rect 20267 21088 20284 21105
rect 20323 21099 20340 21116
rect 20377 21083 20394 21100
rect 20428 21088 20445 21105
rect 23589 21088 23606 21105
rect 25820 21088 25837 21105
rect 25981 21088 25998 21105
rect 7282 21054 7299 21071
rect 9536 21054 9553 21071
rect 18322 21054 18339 21071
rect 23428 21054 23445 21071
rect 4798 21020 4815 21037
rect 20116 20986 20133 21003
rect 24463 20986 24480 21003
rect 26855 20986 26872 21003
rect 4177 20884 4194 20901
rect 6569 20884 6586 20901
rect 8639 20884 8656 20901
rect 20047 20884 20064 20901
rect 7604 20816 7621 20833
rect 10824 20816 10841 20833
rect 13492 20816 13509 20833
rect 19012 20816 19029 20833
rect 22508 20816 22525 20833
rect 24670 20816 24687 20833
rect 27982 20816 27999 20833
rect 3142 20782 3159 20799
rect 5534 20782 5551 20799
rect 7803 20782 7820 20799
rect 10979 20782 10996 20799
rect 11023 20782 11040 20799
rect 11859 20782 11876 20799
rect 13691 20782 13708 20799
rect 19173 20782 19190 20799
rect 21220 20782 21237 20799
rect 22646 20782 22663 20799
rect 24765 20782 24782 20799
rect 28137 20782 28154 20799
rect 28181 20782 28198 20799
rect 3302 20748 3319 20765
rect 3353 20748 3370 20765
rect 5694 20748 5711 20765
rect 5745 20748 5762 20765
rect 7764 20748 7781 20765
rect 13652 20748 13669 20765
rect 19223 20748 19240 20765
rect 21381 20748 21398 20765
rect 21431 20748 21448 20765
rect 22692 20748 22709 20765
rect 22876 20748 22893 20765
rect 24578 20748 24595 20765
rect 24670 20748 24687 20765
rect 24716 20748 24733 20765
rect 14527 20714 14544 20731
rect 22255 20714 22272 20731
rect 22600 20714 22617 20731
rect 29017 20714 29034 20731
rect 4821 20612 4838 20629
rect 7926 20612 7943 20629
rect 15516 20612 15533 20629
rect 24555 20612 24572 20629
rect 3985 20578 4002 20595
rect 15424 20578 15441 20595
rect 21293 20578 21310 20595
rect 22600 20578 22617 20595
rect 23731 20578 23748 20595
rect 25743 20578 25760 20595
rect 28280 20578 28297 20595
rect 29155 20578 29172 20595
rect 3786 20544 3803 20561
rect 3941 20544 3958 20561
rect 6517 20544 6534 20561
rect 6561 20544 6578 20561
rect 7397 20544 7414 20561
rect 7650 20544 7667 20561
rect 7742 20544 7759 20561
rect 7788 20544 7805 20561
rect 7834 20544 7851 20561
rect 11715 20544 11732 20561
rect 11759 20544 11776 20561
rect 14780 20544 14797 20561
rect 14872 20544 14889 20561
rect 15286 20544 15303 20561
rect 15332 20544 15349 20561
rect 15378 20544 15395 20561
rect 21243 20544 21260 20561
rect 22692 20544 22709 20561
rect 22738 20544 22755 20561
rect 22802 20544 22819 20561
rect 23675 20544 23692 20561
rect 25699 20544 25716 20561
rect 26832 20544 26849 20561
rect 26924 20544 26941 20561
rect 28319 20544 28336 20561
rect 29408 20544 29425 20561
rect 29465 20544 29482 20561
rect 29559 20544 29576 20561
rect 29621 20544 29638 20561
rect 29669 20547 29686 20564
rect 29720 20544 29737 20561
rect 6362 20510 6379 20527
rect 11560 20510 11577 20527
rect 14826 20510 14843 20527
rect 21082 20510 21099 20527
rect 22117 20510 22134 20527
rect 23520 20510 23537 20527
rect 25544 20510 25561 20527
rect 28120 20510 28137 20527
rect 22600 20476 22617 20493
rect 26878 20476 26895 20493
rect 12595 20442 12612 20459
rect 26579 20442 26596 20459
rect 29408 20442 29425 20459
rect 6385 20340 6402 20357
rect 14228 20340 14245 20357
rect 17264 20340 17281 20357
rect 26740 20340 26757 20357
rect 29017 20340 29034 20357
rect 11422 20272 11439 20289
rect 12940 20272 12957 20289
rect 15976 20272 15993 20289
rect 19518 20272 19535 20289
rect 5350 20238 5367 20255
rect 5511 20238 5528 20255
rect 11621 20238 11638 20255
rect 13095 20238 13112 20255
rect 13975 20238 13992 20255
rect 14228 20238 14245 20255
rect 14305 20238 14322 20255
rect 14379 20236 14396 20253
rect 14427 20238 14444 20255
rect 14489 20238 14506 20255
rect 14540 20238 14557 20255
rect 16175 20238 16192 20255
rect 17264 20238 17281 20255
rect 17321 20238 17338 20255
rect 17422 20238 17439 20255
rect 17470 20238 17487 20255
rect 17525 20244 17542 20261
rect 17576 20238 17593 20255
rect 26740 20238 26757 20255
rect 26797 20238 26814 20255
rect 26901 20228 26918 20245
rect 26953 20238 26970 20255
rect 27001 20238 27018 20255
rect 27052 20238 27069 20255
rect 27982 20238 27999 20255
rect 28137 20238 28154 20255
rect 5561 20204 5578 20221
rect 11582 20204 11599 20221
rect 13151 20204 13168 20221
rect 16136 20204 16153 20221
rect 17011 20204 17028 20221
rect 19678 20204 19695 20221
rect 19729 20204 19746 20221
rect 28181 20204 28198 20221
rect 12457 20170 12474 20187
rect 20553 20170 20570 20187
rect 13837 20068 13854 20085
rect 6389 20034 6406 20051
rect 9011 20034 9028 20051
rect 10180 20034 10197 20051
rect 12962 20034 12979 20051
rect 13013 20034 13030 20051
rect 15769 20034 15786 20051
rect 17935 20034 17952 20051
rect 20806 20034 20823 20051
rect 23225 20034 23242 20051
rect 25789 20034 25806 20051
rect 6339 20000 6356 20017
rect 7213 20000 7230 20017
rect 8800 20000 8817 20017
rect 8961 20000 8978 20017
rect 10088 20000 10105 20017
rect 10226 20000 10243 20017
rect 10275 20000 10292 20017
rect 11744 20000 11761 20017
rect 11836 20000 11853 20017
rect 11882 20000 11899 20017
rect 11928 20000 11945 20017
rect 12250 20000 12267 20017
rect 12296 20000 12313 20017
rect 12388 20000 12405 20017
rect 12434 20000 12451 20017
rect 12494 20000 12511 20017
rect 15717 20000 15734 20017
rect 16597 20000 16614 20017
rect 17879 20000 17896 20017
rect 19012 20000 19029 20017
rect 19104 20000 19121 20017
rect 20622 20000 20639 20017
rect 20668 20000 20685 20017
rect 20760 20000 20777 20017
rect 20852 20000 20869 20017
rect 23014 20000 23031 20017
rect 23169 20000 23186 20017
rect 24049 20000 24066 20017
rect 24302 20000 24319 20017
rect 24394 20000 24411 20017
rect 24440 20000 24457 20017
rect 24489 20000 24506 20017
rect 25590 20000 25607 20017
rect 25745 20000 25762 20017
rect 26625 20000 26642 20017
rect 6178 19966 6195 19983
rect 9835 19966 9852 19983
rect 12802 19966 12819 19983
rect 15562 19966 15579 19983
rect 17724 19966 17741 19983
rect 18759 19966 18776 19983
rect 12020 19932 12037 19949
rect 12250 19932 12267 19949
rect 10088 19898 10105 19915
rect 19058 19898 19075 19915
rect 20622 19898 20639 19915
rect 24302 19898 24319 19915
rect 9697 19796 9714 19813
rect 11997 19796 12014 19813
rect 14021 19796 14038 19813
rect 17011 19796 17028 19813
rect 5396 19728 5413 19745
rect 8662 19728 8679 19745
rect 10226 19728 10243 19745
rect 10594 19728 10611 19745
rect 10962 19728 10979 19745
rect 19380 19728 19397 19745
rect 5551 19694 5568 19711
rect 8823 19694 8840 19711
rect 10318 19694 10335 19711
rect 10364 19694 10381 19711
rect 11123 19694 11140 19711
rect 12986 19694 13003 19711
rect 13185 19694 13202 19711
rect 15976 19694 15993 19711
rect 16131 19694 16148 19711
rect 21312 19694 21329 19711
rect 21511 19694 21528 19711
rect 5607 19660 5624 19677
rect 8869 19660 8886 19677
rect 11173 19660 11190 19677
rect 13146 19660 13163 19677
rect 16187 19660 16204 19677
rect 19540 19660 19557 19677
rect 19591 19660 19608 19677
rect 21472 19660 21489 19677
rect 6431 19626 6448 19643
rect 20415 19626 20432 19643
rect 22347 19626 22364 19643
rect 20576 19524 20593 19541
rect 22600 19524 22617 19541
rect 24187 19524 24204 19541
rect 3767 19490 3784 19507
rect 7493 19490 7510 19507
rect 8317 19490 8334 19507
rect 20392 19490 20409 19507
rect 20438 19490 20455 19507
rect 21293 19490 21310 19507
rect 23351 19490 23368 19507
rect 3556 19456 3573 19473
rect 3717 19456 3734 19473
rect 4844 19456 4861 19473
rect 4921 19456 4938 19473
rect 5005 19467 5022 19484
rect 5050 19467 5067 19484
rect 5105 19456 5122 19473
rect 5156 19456 5173 19473
rect 7282 19456 7299 19473
rect 7437 19456 7454 19473
rect 8800 19456 8817 19473
rect 8857 19456 8874 19473
rect 8961 19451 8978 19468
rect 9013 19456 9030 19473
rect 9061 19456 9078 19473
rect 9112 19456 9129 19473
rect 20300 19456 20317 19473
rect 20484 19456 20501 19473
rect 21237 19456 21254 19473
rect 22600 19456 22617 19473
rect 22657 19456 22674 19473
rect 22751 19456 22768 19473
rect 22799 19456 22816 19473
rect 22853 19467 22870 19484
rect 22912 19456 22929 19473
rect 23307 19456 23324 19473
rect 4591 19422 4608 19439
rect 21082 19422 21099 19439
rect 22117 19422 22134 19439
rect 23152 19422 23169 19439
rect 8800 19388 8817 19405
rect 4844 19354 4861 19371
rect 4177 19252 4194 19269
rect 6868 19252 6885 19269
rect 8455 19252 8472 19269
rect 19955 19252 19972 19269
rect 22485 19252 22502 19269
rect 27246 19218 27263 19235
rect 5534 19184 5551 19201
rect 7420 19184 7437 19201
rect 18920 19184 18937 19201
rect 27384 19184 27401 19201
rect 3142 19150 3159 19167
rect 3303 19150 3320 19167
rect 6960 19150 6977 19167
rect 7619 19150 7636 19167
rect 19119 19150 19136 19167
rect 21450 19150 21467 19167
rect 21649 19150 21666 19167
rect 24394 19150 24411 19167
rect 24593 19150 24610 19167
rect 27200 19150 27217 19167
rect 3353 19116 3370 19133
rect 5694 19116 5711 19133
rect 5745 19116 5762 19133
rect 6822 19116 6839 19133
rect 6914 19116 6931 19133
rect 7580 19116 7597 19133
rect 19080 19116 19097 19133
rect 21610 19116 21627 19133
rect 24554 19116 24571 19133
rect 6569 19082 6586 19099
rect 25429 19082 25446 19099
rect 27246 19082 27263 19099
rect 27292 19082 27309 19099
rect 6454 18980 6471 18997
rect 8317 18980 8334 18997
rect 24394 18980 24411 18997
rect 24762 18980 24779 18997
rect 24808 18980 24825 18997
rect 3629 18946 3646 18963
rect 4706 18946 4723 18963
rect 6500 18946 6517 18963
rect 6546 18946 6563 18963
rect 7493 18946 7510 18963
rect 12047 18946 12064 18963
rect 14480 18946 14497 18963
rect 14531 18946 14548 18963
rect 17889 18946 17906 18963
rect 23133 18946 23150 18963
rect 25498 18946 25515 18963
rect 26491 18946 26508 18963
rect 28423 18946 28440 18963
rect 3418 18912 3435 18929
rect 3573 18912 3590 18929
rect 4798 18912 4815 18929
rect 4844 18912 4861 18929
rect 6362 18912 6379 18929
rect 6408 18912 6425 18929
rect 6592 18912 6609 18929
rect 7282 18912 7299 18929
rect 7437 18912 7454 18929
rect 11991 18912 12008 18929
rect 15355 18912 15372 18929
rect 15608 18912 15625 18929
rect 15700 18912 15717 18929
rect 15746 18912 15763 18929
rect 15795 18912 15812 18929
rect 17678 18912 17695 18929
rect 17839 18912 17856 18929
rect 23083 18912 23100 18929
rect 24302 18912 24319 18929
rect 24348 18912 24365 18929
rect 24486 18912 24503 18929
rect 24716 18912 24733 18929
rect 25360 18912 25377 18929
rect 25452 18912 25469 18929
rect 25547 18907 25564 18924
rect 26435 18912 26452 18929
rect 28212 18912 28229 18929
rect 28367 18912 28384 18929
rect 29247 18912 29264 18929
rect 29500 18912 29517 18929
rect 29592 18912 29609 18929
rect 29638 18912 29655 18929
rect 29687 18912 29704 18929
rect 11836 18878 11853 18895
rect 14320 18878 14337 18895
rect 22922 18878 22939 18895
rect 24900 18878 24917 18895
rect 25406 18878 25423 18895
rect 26280 18878 26297 18895
rect 29546 18878 29563 18895
rect 4844 18844 4861 18861
rect 24210 18844 24227 18861
rect 4453 18810 4470 18827
rect 12871 18810 12888 18827
rect 15608 18810 15625 18827
rect 18713 18810 18730 18827
rect 23957 18810 23974 18827
rect 24762 18810 24779 18827
rect 27315 18810 27332 18827
rect 4660 18708 4677 18725
rect 10870 18708 10887 18725
rect 15217 18708 15234 18725
rect 25291 18708 25308 18725
rect 27384 18708 27401 18725
rect 20530 18674 20547 18691
rect 13032 18640 13049 18657
rect 26188 18640 26205 18657
rect 27982 18640 27999 18657
rect 4862 18606 4879 18623
rect 5258 18606 5275 18623
rect 5419 18606 5436 18623
rect 8294 18606 8311 18623
rect 8455 18606 8472 18623
rect 10962 18606 10979 18623
rect 11057 18606 11074 18623
rect 11422 18606 11439 18623
rect 13078 18606 13095 18623
rect 13127 18606 13144 18623
rect 14182 18606 14199 18623
rect 14337 18606 14354 18623
rect 15700 18606 15717 18623
rect 15884 18606 15901 18623
rect 16160 18606 16177 18623
rect 16359 18606 16376 18623
rect 19242 18606 19259 18623
rect 19397 18606 19414 18623
rect 20717 18606 20734 18623
rect 21220 18606 21237 18623
rect 21404 18606 21421 18623
rect 21956 18606 21973 18623
rect 22033 18606 22050 18623
rect 22114 18606 22131 18623
rect 22169 18606 22186 18623
rect 22217 18604 22234 18621
rect 22268 18606 22285 18623
rect 24256 18606 24273 18623
rect 26096 18606 26113 18623
rect 27476 18606 27493 18623
rect 27571 18606 27588 18623
rect 28137 18606 28154 18623
rect 4660 18572 4677 18589
rect 4752 18572 4769 18589
rect 4798 18572 4815 18589
rect 5469 18572 5486 18589
rect 8505 18572 8522 18589
rect 10870 18572 10887 18589
rect 11008 18572 11025 18589
rect 11582 18572 11599 18589
rect 11633 18572 11650 18589
rect 12457 18572 12474 18589
rect 12940 18572 12957 18589
rect 13032 18572 13049 18589
rect 14393 18572 14410 18589
rect 16320 18572 16337 18589
rect 19453 18572 19470 18589
rect 20277 18572 20294 18589
rect 20530 18572 20547 18589
rect 20622 18572 20639 18589
rect 20668 18572 20685 18589
rect 24416 18572 24433 18589
rect 24467 18572 24484 18589
rect 26234 18572 26251 18589
rect 26280 18572 26297 18589
rect 27384 18572 27401 18589
rect 27522 18572 27539 18589
rect 28189 18572 28206 18589
rect 6293 18538 6310 18555
rect 9329 18538 9346 18555
rect 15746 18538 15763 18555
rect 15792 18538 15809 18555
rect 15838 18538 15855 18555
rect 17195 18538 17212 18555
rect 21266 18538 21283 18555
rect 21312 18538 21329 18555
rect 21358 18538 21375 18555
rect 21956 18538 21973 18555
rect 29017 18538 29034 18555
rect 4361 18436 4378 18453
rect 6224 18436 6241 18453
rect 6270 18436 6287 18453
rect 11031 18436 11048 18453
rect 16528 18436 16545 18453
rect 19357 18436 19374 18453
rect 21795 18436 21812 18453
rect 24049 18436 24066 18453
rect 29431 18436 29448 18453
rect 3537 18402 3554 18419
rect 6895 18402 6912 18419
rect 10207 18402 10224 18419
rect 13009 18402 13026 18419
rect 15354 18402 15371 18419
rect 16229 18402 16246 18419
rect 17080 18402 17097 18419
rect 18533 18402 18550 18419
rect 23221 18402 23238 18419
rect 24302 18402 24319 18419
rect 24440 18402 24457 18419
rect 28556 18402 28573 18419
rect 28607 18402 28624 18419
rect 3326 18368 3343 18385
rect 3487 18368 3504 18385
rect 6845 18368 6862 18385
rect 9352 18368 9369 18385
rect 9409 18368 9426 18385
rect 9503 18368 9520 18385
rect 9551 18379 9568 18396
rect 9613 18368 9630 18385
rect 9664 18368 9681 18385
rect 10151 18368 10168 18385
rect 12963 18368 12980 18385
rect 15393 18368 15410 18385
rect 16482 18368 16499 18385
rect 16574 18368 16591 18385
rect 17172 18368 17189 18385
rect 17218 18368 17235 18385
rect 17267 18368 17284 18385
rect 18477 18368 18494 18385
rect 20915 18368 20932 18385
rect 20959 18368 20976 18385
rect 23169 18368 23186 18385
rect 24394 18368 24411 18385
rect 24489 18368 24506 18385
rect 6316 18334 6333 18351
rect 6684 18334 6701 18351
rect 9996 18334 10013 18351
rect 12802 18334 12819 18351
rect 15194 18334 15211 18351
rect 17080 18334 17097 18351
rect 18322 18334 18339 18351
rect 20760 18334 20777 18351
rect 23014 18334 23031 18351
rect 24348 18334 24365 18351
rect 28396 18334 28413 18351
rect 9352 18300 9369 18317
rect 6040 18266 6057 18283
rect 7719 18266 7736 18283
rect 13837 18266 13854 18283
rect 4177 18164 4194 18181
rect 6040 18164 6057 18181
rect 7420 18164 7437 18181
rect 9467 18164 9484 18181
rect 11215 18164 11232 18181
rect 17241 18164 17258 18181
rect 22255 18164 22272 18181
rect 5166 18096 5183 18113
rect 5304 18096 5321 18113
rect 14435 18096 14452 18113
rect 3142 18062 3159 18079
rect 3297 18062 3314 18079
rect 6684 18062 6701 18079
rect 6868 18062 6885 18079
rect 7420 18062 7437 18079
rect 7466 18062 7483 18079
rect 7650 18062 7667 18079
rect 8432 18062 8449 18079
rect 8587 18062 8604 18079
rect 10180 18062 10197 18079
rect 10335 18062 10352 18079
rect 13400 18062 13417 18079
rect 13561 18062 13578 18079
rect 14688 18062 14705 18079
rect 14765 18062 14782 18079
rect 14839 18062 14856 18079
rect 14887 18062 14904 18079
rect 14949 18068 14966 18085
rect 15000 18062 15017 18079
rect 16206 18062 16223 18079
rect 21220 18062 21237 18079
rect 3353 18028 3370 18045
rect 6776 18028 6793 18045
rect 6822 18028 6839 18045
rect 7558 18028 7575 18045
rect 7604 18028 7621 18045
rect 8631 18028 8648 18045
rect 10391 18028 10408 18045
rect 13611 18028 13628 18045
rect 16366 18028 16383 18045
rect 16417 18028 16434 18045
rect 21380 18028 21397 18045
rect 21431 18028 21448 18045
rect 6960 17994 6977 18011
rect 14918 17994 14935 18011
rect 13837 17892 13854 17909
rect 22117 17892 22134 17909
rect 24256 17892 24273 17909
rect 6844 17858 6861 17875
rect 6895 17858 6912 17875
rect 13013 17858 13030 17875
rect 21293 17858 21310 17875
rect 22949 17858 22966 17875
rect 26445 17858 26462 17875
rect 6684 17824 6701 17841
rect 12802 17824 12819 17841
rect 12957 17824 12974 17841
rect 18782 17824 18799 17841
rect 18874 17824 18891 17841
rect 21243 17824 21260 17841
rect 22893 17824 22910 17841
rect 24026 17824 24043 17841
rect 24083 17824 24100 17841
rect 24177 17824 24194 17841
rect 24239 17824 24256 17841
rect 24287 17824 24304 17841
rect 24338 17824 24355 17841
rect 26389 17824 26406 17841
rect 7719 17790 7736 17807
rect 21082 17790 21099 17807
rect 22738 17790 22755 17807
rect 23773 17790 23790 17807
rect 26234 17790 26251 17807
rect 18828 17722 18845 17739
rect 27269 17722 27286 17739
rect 4660 17620 4677 17637
rect 6661 17620 6678 17637
rect 9283 17620 9300 17637
rect 18782 17620 18799 17637
rect 23497 17620 23514 17637
rect 25774 17620 25791 17637
rect 3142 17552 3159 17569
rect 8248 17552 8265 17569
rect 22462 17552 22479 17569
rect 4752 17518 4769 17535
rect 4862 17518 4879 17535
rect 5626 17518 5643 17535
rect 5781 17518 5798 17535
rect 8409 17518 8426 17535
rect 18782 17518 18799 17535
rect 18839 17518 18856 17535
rect 18933 17518 18950 17535
rect 18995 17508 19012 17525
rect 19043 17516 19060 17533
rect 19094 17518 19111 17535
rect 22623 17518 22640 17535
rect 24486 17518 24503 17535
rect 24647 17518 24664 17535
rect 25774 17518 25791 17535
rect 25851 17518 25868 17535
rect 25932 17518 25949 17535
rect 25980 17508 25997 17525
rect 26035 17518 26052 17535
rect 26086 17518 26103 17535
rect 27982 17518 27999 17535
rect 3302 17484 3319 17501
rect 3353 17484 3370 17501
rect 4177 17484 4194 17501
rect 4660 17484 4677 17501
rect 4798 17484 4815 17501
rect 5837 17484 5854 17501
rect 8459 17484 8476 17501
rect 22673 17484 22690 17501
rect 24693 17484 24710 17501
rect 25521 17484 25538 17501
rect 28142 17484 28159 17501
rect 28193 17484 28210 17501
rect 29017 17450 29034 17467
rect 4637 17348 4654 17365
rect 18759 17348 18776 17365
rect 26395 17348 26412 17365
rect 3813 17314 3830 17331
rect 7447 17314 7464 17331
rect 12829 17314 12846 17331
rect 14887 17314 14904 17331
rect 17935 17314 17952 17331
rect 20465 17314 20482 17331
rect 23179 17314 23196 17331
rect 25571 17314 25588 17331
rect 28423 17314 28440 17331
rect 29500 17314 29517 17331
rect 3763 17280 3780 17297
rect 7236 17280 7253 17297
rect 7397 17280 7414 17297
rect 12779 17280 12796 17297
rect 14843 17280 14860 17297
rect 17724 17280 17741 17297
rect 17879 17280 17896 17297
rect 20409 17280 20426 17297
rect 23123 17280 23140 17297
rect 25521 17280 25538 17297
rect 27108 17280 27125 17297
rect 27165 17280 27182 17297
rect 27266 17280 27283 17297
rect 27321 17291 27338 17308
rect 27369 17280 27386 17297
rect 27420 17280 27437 17297
rect 28367 17280 28384 17297
rect 29592 17280 29609 17297
rect 29638 17280 29655 17297
rect 29702 17280 29719 17297
rect 3602 17246 3619 17263
rect 12618 17246 12635 17263
rect 14688 17246 14705 17263
rect 20254 17246 20271 17263
rect 22968 17246 22985 17263
rect 25360 17246 25377 17263
rect 28212 17246 28229 17263
rect 29247 17246 29264 17263
rect 24003 17212 24020 17229
rect 8271 17178 8288 17195
rect 13653 17178 13670 17195
rect 15723 17178 15740 17195
rect 21289 17178 21306 17195
rect 27108 17178 27125 17195
rect 29500 17178 29517 17195
rect 6523 17076 6540 17093
rect 25567 17076 25584 17093
rect 27775 17076 27792 17093
rect 5488 17008 5505 17025
rect 8662 17008 8679 17025
rect 10962 17008 10979 17025
rect 11997 17008 12014 17025
rect 12940 17008 12957 17025
rect 14780 17008 14797 17025
rect 21220 17008 21237 17025
rect 24532 17008 24549 17025
rect 28626 17008 28643 17025
rect 5649 16974 5666 16991
rect 8823 16974 8840 16991
rect 12250 16974 12267 16991
rect 12342 16974 12359 16991
rect 14734 16974 14751 16991
rect 14844 16974 14861 16991
rect 15148 16974 15165 16991
rect 15240 16974 15257 16991
rect 15792 16974 15809 16991
rect 17080 16974 17097 16991
rect 17172 16974 17189 16991
rect 21381 16974 21398 16991
rect 24687 16974 24704 16991
rect 26740 16974 26757 16991
rect 28718 16974 28735 16991
rect 5699 16940 5716 16957
rect 8869 16940 8886 16957
rect 11122 16940 11139 16957
rect 11173 16940 11190 16957
rect 13100 16940 13117 16957
rect 13151 16940 13168 16957
rect 14642 16940 14659 16957
rect 14780 16940 14797 16957
rect 15952 16940 15969 16957
rect 16003 16940 16020 16957
rect 21431 16940 21448 16957
rect 24731 16940 24748 16957
rect 26901 16940 26918 16957
rect 26951 16940 26968 16957
rect 28810 16940 28827 16957
rect 28994 16940 29011 16957
rect 9697 16906 9714 16923
rect 12296 16906 12313 16923
rect 13975 16906 13992 16923
rect 15194 16906 15211 16923
rect 16827 16906 16844 16923
rect 17172 16906 17189 16923
rect 22255 16906 22272 16923
rect 28764 16906 28781 16923
rect 13837 16804 13854 16821
rect 14550 16804 14567 16821
rect 14964 16804 14981 16821
rect 15010 16804 15027 16821
rect 15056 16804 15073 16821
rect 18805 16804 18822 16821
rect 21312 16804 21329 16821
rect 27039 16804 27056 16821
rect 7493 16770 7510 16787
rect 10241 16770 10258 16787
rect 11652 16770 11669 16787
rect 13013 16770 13030 16787
rect 14872 16770 14889 16787
rect 15769 16770 15786 16787
rect 17080 16770 17097 16787
rect 17981 16770 17998 16787
rect 20235 16770 20252 16787
rect 23175 16770 23192 16787
rect 26211 16770 26228 16787
rect 28556 16770 28573 16787
rect 28607 16770 28624 16787
rect 7443 16736 7460 16753
rect 9536 16736 9553 16753
rect 9628 16736 9645 16753
rect 9674 16736 9691 16753
rect 9720 16736 9737 16753
rect 10042 16736 10059 16753
rect 10197 16736 10214 16753
rect 11077 16736 11094 16753
rect 11560 16736 11577 16753
rect 11698 16736 11715 16753
rect 11747 16736 11764 16753
rect 12020 16736 12037 16753
rect 12112 16736 12129 16753
rect 12802 16736 12819 16753
rect 12957 16736 12974 16753
rect 14320 16736 14337 16753
rect 14377 16736 14394 16753
rect 14471 16736 14488 16753
rect 14533 16731 14550 16748
rect 14581 16736 14598 16753
rect 14632 16736 14649 16753
rect 15723 16736 15740 16753
rect 17172 16736 17189 16753
rect 17218 16736 17235 16753
rect 17267 16731 17284 16748
rect 17770 16736 17787 16753
rect 17931 16736 17948 16753
rect 20179 16736 20196 16753
rect 21312 16736 21329 16753
rect 21369 16736 21386 16753
rect 21463 16736 21480 16753
rect 21525 16731 21542 16748
rect 21573 16736 21590 16753
rect 21624 16736 21641 16753
rect 23123 16736 23140 16753
rect 26165 16736 26182 16753
rect 28396 16736 28413 16753
rect 7282 16702 7299 16719
rect 11606 16702 11623 16719
rect 15562 16702 15579 16719
rect 16597 16702 16614 16719
rect 20024 16702 20041 16719
rect 21059 16702 21076 16719
rect 22968 16702 22985 16719
rect 26004 16702 26021 16719
rect 8317 16634 8334 16651
rect 9812 16634 9829 16651
rect 12066 16634 12083 16651
rect 15148 16634 15165 16651
rect 17080 16634 17097 16651
rect 24003 16634 24020 16651
rect 29431 16634 29448 16651
rect 9697 16532 9714 16549
rect 11629 16532 11646 16549
rect 14849 16532 14866 16549
rect 16965 16532 16982 16549
rect 23980 16532 23997 16549
rect 29500 16532 29517 16549
rect 4660 16498 4677 16515
rect 10180 16498 10197 16515
rect 7650 16464 7667 16481
rect 10594 16464 10611 16481
rect 13814 16464 13831 16481
rect 15930 16464 15947 16481
rect 4660 16430 4677 16447
rect 4737 16430 4754 16447
rect 4811 16430 4828 16447
rect 4859 16430 4876 16447
rect 4921 16430 4938 16447
rect 4972 16428 4989 16445
rect 5718 16430 5735 16447
rect 7420 16430 7437 16447
rect 8018 16430 8035 16447
rect 8662 16430 8679 16447
rect 8861 16430 8878 16447
rect 10180 16430 10197 16447
rect 10318 16430 10335 16447
rect 10793 16430 10810 16447
rect 13969 16430 13986 16447
rect 16085 16430 16102 16447
rect 16129 16430 16146 16447
rect 17218 16430 17235 16447
rect 17310 16430 17327 16447
rect 24072 16430 24089 16447
rect 24118 16430 24135 16447
rect 24182 16430 24199 16447
rect 29592 16430 29609 16447
rect 29638 16430 29655 16447
rect 29687 16430 29704 16447
rect 5878 16396 5895 16413
rect 5929 16396 5946 16413
rect 8822 16396 8839 16413
rect 10754 16396 10771 16413
rect 14025 16396 14042 16413
rect 23980 16396 23997 16413
rect 29500 16396 29517 16413
rect 6753 16362 6770 16379
rect 10272 16362 10289 16379
rect 17264 16362 17281 16379
rect 4269 16260 4286 16277
rect 6408 16260 6425 16277
rect 6730 16260 6747 16277
rect 9835 16260 9852 16277
rect 13745 16260 13762 16277
rect 23865 16260 23882 16277
rect 29339 16260 29356 16277
rect 4729 16226 4746 16243
rect 6224 16226 6241 16243
rect 6638 16226 6655 16243
rect 7447 16226 7464 16243
rect 9011 16226 9028 16243
rect 12921 16226 12938 16243
rect 20967 16226 20984 16243
rect 23041 16226 23058 16243
rect 26119 16226 26136 16243
rect 28511 16226 28528 16243
rect 3234 16192 3251 16209
rect 3389 16192 3406 16209
rect 3433 16192 3450 16209
rect 4522 16192 4539 16209
rect 4683 16192 4700 16209
rect 5557 16192 5574 16209
rect 6132 16192 6149 16209
rect 6270 16192 6287 16209
rect 6316 16192 6333 16209
rect 6776 16192 6793 16209
rect 7236 16192 7253 16209
rect 7397 16192 7414 16209
rect 8800 16192 8817 16209
rect 8955 16192 8972 16209
rect 12710 16192 12727 16209
rect 12865 16192 12882 16209
rect 20921 16192 20938 16209
rect 22985 16192 23002 16209
rect 26067 16192 26084 16209
rect 28459 16192 28476 16209
rect 20760 16158 20777 16175
rect 22830 16158 22847 16175
rect 25912 16158 25929 16175
rect 28304 16158 28321 16175
rect 6638 16090 6655 16107
rect 8271 16090 8288 16107
rect 21795 16090 21812 16107
rect 26947 16090 26964 16107
rect 4177 15988 4194 16005
rect 6201 15988 6218 16005
rect 3142 15920 3159 15937
rect 26740 15920 26757 15937
rect 3303 15886 3320 15903
rect 5166 15886 5183 15903
rect 8110 15886 8127 15903
rect 8187 15886 8204 15903
rect 8261 15884 8278 15901
rect 8317 15876 8334 15893
rect 8371 15886 8388 15903
rect 8422 15886 8439 15903
rect 10778 15886 10795 15903
rect 10977 15886 10994 15903
rect 24348 15886 24365 15903
rect 25636 15886 25653 15903
rect 25713 15886 25730 15903
rect 25794 15886 25811 15903
rect 25849 15876 25866 15893
rect 25897 15876 25914 15893
rect 25948 15886 25965 15903
rect 28718 15886 28735 15903
rect 28810 15886 28827 15903
rect 28948 15886 28965 15903
rect 3353 15852 3370 15869
rect 5326 15852 5343 15869
rect 5377 15852 5394 15869
rect 10938 15852 10955 15869
rect 24508 15852 24525 15869
rect 24559 15852 24576 15869
rect 25383 15852 25400 15869
rect 26901 15852 26918 15869
rect 26951 15852 26968 15869
rect 28764 15852 28781 15869
rect 8110 15818 8127 15835
rect 11813 15818 11830 15835
rect 25866 15818 25883 15835
rect 27775 15818 27792 15835
rect 4499 15716 4516 15733
rect 26395 15716 26412 15733
rect 27384 15716 27401 15733
rect 3675 15682 3692 15699
rect 9425 15682 9442 15699
rect 12691 15682 12708 15699
rect 18533 15682 18550 15699
rect 20281 15682 20298 15699
rect 25571 15682 25588 15699
rect 3625 15648 3642 15665
rect 9369 15648 9386 15665
rect 12635 15648 12652 15665
rect 15487 15648 15504 15665
rect 15531 15648 15548 15665
rect 18483 15648 18500 15665
rect 20231 15648 20248 15665
rect 21105 15648 21122 15665
rect 21588 15648 21605 15665
rect 21645 15648 21662 15665
rect 21739 15648 21756 15665
rect 21795 15648 21812 15665
rect 21849 15659 21866 15676
rect 21900 15648 21917 15665
rect 25360 15648 25377 15665
rect 25521 15648 25538 15665
rect 27154 15648 27171 15665
rect 27211 15648 27228 15665
rect 27305 15651 27322 15668
rect 27353 15648 27370 15665
rect 27415 15648 27432 15665
rect 27466 15648 27483 15665
rect 3464 15614 3481 15631
rect 9214 15614 9231 15631
rect 12480 15614 12497 15631
rect 15332 15614 15349 15631
rect 18322 15614 18339 15631
rect 20070 15614 20087 15631
rect 10249 15546 10266 15563
rect 13515 15546 13532 15563
rect 16367 15546 16384 15563
rect 19357 15546 19374 15563
rect 21588 15546 21605 15563
rect 17977 15444 17994 15461
rect 25291 15444 25308 15461
rect 27775 15444 27792 15461
rect 5580 15376 5597 15393
rect 10870 15376 10887 15393
rect 15930 15376 15947 15393
rect 16252 15376 16269 15393
rect 18460 15376 18477 15393
rect 20070 15376 20087 15393
rect 22830 15376 22847 15393
rect 24256 15376 24273 15393
rect 26740 15376 26757 15393
rect 5741 15342 5758 15359
rect 7834 15342 7851 15359
rect 7995 15342 8012 15359
rect 11025 15342 11042 15359
rect 13814 15342 13831 15359
rect 13969 15342 13986 15359
rect 15884 15342 15901 15359
rect 15979 15342 15996 15359
rect 16439 15342 16456 15359
rect 16942 15342 16959 15359
rect 18621 15342 18638 15359
rect 19495 15342 19512 15359
rect 20116 15342 20133 15359
rect 20165 15342 20182 15359
rect 22738 15342 22755 15359
rect 22922 15342 22939 15359
rect 24411 15342 24428 15359
rect 26895 15342 26912 15359
rect 5791 15308 5808 15325
rect 8045 15308 8062 15325
rect 11081 15308 11098 15325
rect 14025 15308 14042 15325
rect 15792 15308 15809 15325
rect 15930 15308 15947 15325
rect 16252 15308 16269 15325
rect 16344 15308 16361 15325
rect 16390 15308 16407 15325
rect 17102 15308 17119 15325
rect 17153 15308 17170 15325
rect 18671 15308 18688 15325
rect 19978 15308 19995 15325
rect 20070 15308 20087 15325
rect 22784 15308 22801 15325
rect 24455 15308 24472 15325
rect 26951 15308 26968 15325
rect 6615 15274 6632 15291
rect 8869 15274 8886 15291
rect 11905 15274 11922 15291
rect 14849 15274 14866 15291
rect 22876 15274 22893 15291
rect 6454 15172 6471 15189
rect 16413 15172 16430 15189
rect 21565 15172 21582 15189
rect 3767 15138 3784 15155
rect 4936 15138 4953 15155
rect 6868 15138 6885 15155
rect 7442 15138 7459 15155
rect 10249 15138 10266 15155
rect 11077 15138 11094 15155
rect 12962 15138 12979 15155
rect 13013 15138 13030 15155
rect 13837 15138 13854 15155
rect 15589 15138 15606 15155
rect 20741 15138 20758 15155
rect 28557 15138 28574 15155
rect 3711 15104 3728 15121
rect 4844 15104 4861 15121
rect 4982 15104 4999 15121
rect 5028 15104 5045 15121
rect 6362 15104 6379 15121
rect 6408 15104 6425 15121
rect 6546 15104 6563 15121
rect 6776 15104 6793 15121
rect 6914 15104 6931 15121
rect 6960 15104 6977 15121
rect 7481 15104 7498 15121
rect 8800 15104 8817 15121
rect 8857 15104 8874 15121
rect 8951 15104 8968 15121
rect 9013 15104 9030 15121
rect 9061 15115 9078 15132
rect 9112 15104 9129 15121
rect 10203 15104 10220 15121
rect 11698 15104 11715 15121
rect 11755 15104 11772 15121
rect 11849 15104 11866 15121
rect 11911 15104 11928 15121
rect 11959 15104 11976 15121
rect 12010 15107 12027 15124
rect 14458 15104 14475 15121
rect 14515 15104 14532 15121
rect 14609 15107 14626 15124
rect 14657 15099 14674 15116
rect 14719 15099 14736 15116
rect 14770 15104 14787 15121
rect 15533 15104 15550 15121
rect 18506 15104 18523 15121
rect 18920 15104 18937 15121
rect 20530 15104 20547 15121
rect 20691 15104 20708 15121
rect 28350 15104 28367 15121
rect 28505 15104 28522 15121
rect 3556 15070 3573 15087
rect 7282 15070 7299 15087
rect 8317 15070 8334 15087
rect 10042 15070 10059 15087
rect 12802 15070 12819 15087
rect 15378 15070 15395 15087
rect 18736 15070 18753 15087
rect 4591 15002 4608 15019
rect 5120 15002 5137 15019
rect 6408 15002 6425 15019
rect 7052 15002 7069 15019
rect 8800 15002 8817 15019
rect 11698 15002 11715 15019
rect 14458 15002 14475 15019
rect 29385 15002 29402 15019
rect 4177 14900 4194 14917
rect 7420 14900 7437 14917
rect 15217 14900 15234 14917
rect 16114 14900 16131 14917
rect 3142 14832 3159 14849
rect 6937 14832 6954 14849
rect 11422 14832 11439 14849
rect 14182 14832 14199 14849
rect 16160 14832 16177 14849
rect 24624 14832 24641 14849
rect 4752 14798 4769 14815
rect 4798 14798 4815 14815
rect 4982 14798 4999 14815
rect 5902 14798 5919 14815
rect 6057 14798 6074 14815
rect 7420 14798 7437 14815
rect 7466 14798 7483 14815
rect 7604 14798 7621 14815
rect 7650 14798 7667 14815
rect 8662 14798 8679 14815
rect 8823 14798 8840 14815
rect 10180 14798 10197 14815
rect 10237 14798 10254 14815
rect 10341 14788 10358 14805
rect 10393 14798 10410 14815
rect 10441 14804 10458 14821
rect 10492 14798 10509 14815
rect 11583 14798 11600 14815
rect 13400 14798 13417 14815
rect 13457 14798 13474 14815
rect 13551 14796 13568 14813
rect 13599 14804 13616 14821
rect 13661 14798 13678 14815
rect 13712 14798 13729 14815
rect 15976 14798 15993 14815
rect 24779 14798 24796 14815
rect 3302 14764 3319 14781
rect 3353 14764 3370 14781
rect 4890 14764 4907 14781
rect 4936 14764 4953 14781
rect 6113 14764 6130 14781
rect 7558 14764 7575 14781
rect 8869 14764 8886 14781
rect 9697 14764 9714 14781
rect 11633 14764 11650 14781
rect 12457 14764 12474 14781
rect 14342 14764 14359 14781
rect 14393 14764 14410 14781
rect 16022 14764 16039 14781
rect 24831 14764 24848 14781
rect 4844 14730 4861 14747
rect 10180 14730 10197 14747
rect 13630 14730 13647 14747
rect 16068 14730 16085 14747
rect 25659 14730 25676 14747
rect 4821 14628 4838 14645
rect 7719 14628 7736 14645
rect 13423 14628 13440 14645
rect 3985 14594 4002 14611
rect 6895 14594 6912 14611
rect 9333 14594 9350 14611
rect 12599 14594 12616 14611
rect 15405 14594 15422 14611
rect 26399 14594 26416 14611
rect 3941 14560 3958 14577
rect 6839 14560 6856 14577
rect 9277 14560 9294 14577
rect 12388 14560 12405 14577
rect 12543 14560 12560 14577
rect 15349 14560 15366 14577
rect 26349 14560 26366 14577
rect 29362 14560 29379 14577
rect 29454 14560 29471 14577
rect 3786 14526 3803 14543
rect 6684 14526 6701 14543
rect 9122 14526 9139 14543
rect 15194 14526 15211 14543
rect 26188 14526 26205 14543
rect 10157 14458 10174 14475
rect 16229 14458 16246 14475
rect 27223 14458 27240 14475
rect 29408 14458 29425 14475
rect 4177 14356 4194 14373
rect 6799 14356 6816 14373
rect 8685 14356 8702 14373
rect 14297 14356 14314 14373
rect 22876 14322 22893 14339
rect 3142 14288 3159 14305
rect 5764 14288 5781 14305
rect 7650 14288 7667 14305
rect 11905 14288 11922 14305
rect 17310 14288 17327 14305
rect 17770 14288 17787 14305
rect 21220 14288 21237 14305
rect 21358 14288 21375 14305
rect 24348 14288 24365 14305
rect 25383 14288 25400 14305
rect 3297 14254 3314 14271
rect 5925 14254 5942 14271
rect 7805 14254 7822 14271
rect 7849 14254 7866 14271
rect 10870 14254 10887 14271
rect 11031 14254 11048 14271
rect 12158 14254 12175 14271
rect 12204 14254 12221 14271
rect 12342 14254 12359 14271
rect 12388 14254 12405 14271
rect 13262 14254 13279 14271
rect 13461 14254 13478 14271
rect 17678 14254 17695 14271
rect 17862 14254 17879 14271
rect 19518 14254 19535 14271
rect 19932 14254 19949 14271
rect 21266 14254 21283 14271
rect 22876 14254 22893 14271
rect 23014 14254 23031 14271
rect 25636 14254 25653 14271
rect 25693 14254 25710 14271
rect 25787 14254 25804 14271
rect 25835 14254 25852 14271
rect 25890 14252 25907 14269
rect 25948 14254 25965 14271
rect 27706 14254 27723 14271
rect 27861 14254 27878 14271
rect 3353 14220 3370 14237
rect 5975 14220 5992 14237
rect 11081 14220 11098 14237
rect 12296 14220 12313 14237
rect 13422 14220 13439 14237
rect 19702 14220 19719 14237
rect 22968 14220 22985 14237
rect 24508 14220 24525 14237
rect 24559 14220 24576 14237
rect 27917 14220 27934 14237
rect 12250 14186 12267 14203
rect 17402 14186 17419 14203
rect 17724 14186 17741 14203
rect 17816 14186 17833 14203
rect 19518 14186 19535 14203
rect 21358 14186 21375 14203
rect 25866 14186 25883 14203
rect 28741 14186 28758 14203
rect 17770 14084 17787 14101
rect 21450 14084 21467 14101
rect 4733 14050 4750 14067
rect 9720 14050 9737 14067
rect 26169 14050 26186 14067
rect 28331 14050 28348 14067
rect 4683 14016 4700 14033
rect 6086 14016 6103 14033
rect 6133 14016 6150 14033
rect 6224 14016 6241 14033
rect 6270 14016 6287 14033
rect 6339 14016 6356 14033
rect 9628 14016 9645 14033
rect 9766 14016 9783 14033
rect 9830 14016 9847 14033
rect 15240 14016 15257 14033
rect 15286 14016 15303 14033
rect 15378 14016 15395 14033
rect 15424 14016 15441 14033
rect 15470 14016 15487 14033
rect 17208 14016 17225 14033
rect 19886 14016 19903 14033
rect 20300 14016 20317 14033
rect 20530 14016 20547 14033
rect 20622 14016 20639 14033
rect 21358 14016 21375 14033
rect 21404 14016 21421 14033
rect 26113 14016 26130 14033
rect 26993 14016 27010 14033
rect 27246 14016 27263 14033
rect 27303 14016 27320 14033
rect 27397 14016 27414 14033
rect 27445 14011 27462 14028
rect 27500 14027 27517 14044
rect 27558 14016 27575 14033
rect 28275 14016 28292 14033
rect 4522 13982 4539 13999
rect 5557 13982 5574 13999
rect 17080 13982 17097 13999
rect 20070 13982 20087 13999
rect 21542 13982 21559 13999
rect 25958 13982 25975 13999
rect 28120 13982 28137 13999
rect 20576 13948 20593 13965
rect 21404 13948 21421 13965
rect 6408 13914 6425 13931
rect 9628 13914 9645 13931
rect 15240 13914 15257 13931
rect 27246 13914 27263 13931
rect 29155 13914 29172 13931
rect 6201 13812 6218 13829
rect 9513 13812 9530 13829
rect 11721 13812 11738 13829
rect 15217 13812 15234 13829
rect 16758 13812 16775 13829
rect 25521 13812 25538 13829
rect 23014 13778 23031 13795
rect 26832 13778 26849 13795
rect 8478 13744 8495 13761
rect 16804 13744 16821 13761
rect 18690 13744 18707 13761
rect 24486 13744 24503 13761
rect 26970 13744 26987 13761
rect 28626 13744 28643 13761
rect 5166 13710 5183 13727
rect 8639 13710 8656 13727
rect 10686 13710 10703 13727
rect 10847 13710 10864 13727
rect 14182 13710 14199 13727
rect 14337 13710 14354 13727
rect 16666 13710 16683 13727
rect 16712 13710 16729 13727
rect 23106 13710 23123 13727
rect 23152 13710 23169 13727
rect 24641 13710 24658 13727
rect 26786 13710 26803 13727
rect 26832 13710 26849 13727
rect 28828 13710 28845 13727
rect 29500 13710 29517 13727
rect 29592 13710 29609 13727
rect 5326 13676 5343 13693
rect 5377 13676 5394 13693
rect 8689 13676 8706 13693
rect 10897 13676 10914 13693
rect 14393 13676 14410 13693
rect 18824 13676 18841 13693
rect 23014 13676 23031 13693
rect 24697 13676 24714 13693
rect 28626 13676 28643 13693
rect 28718 13676 28735 13693
rect 28764 13676 28781 13693
rect 19380 13642 19397 13659
rect 26878 13642 26895 13659
rect 29546 13642 29563 13659
rect 9674 13540 9691 13557
rect 15355 13540 15372 13557
rect 16298 13540 16315 13557
rect 27039 13540 27056 13557
rect 3537 13506 3554 13523
rect 4361 13506 4378 13523
rect 4752 13506 4769 13523
rect 5074 13506 5091 13523
rect 7074 13506 7091 13523
rect 7125 13506 7142 13523
rect 9582 13506 9599 13523
rect 9628 13506 9645 13523
rect 10253 13506 10270 13523
rect 13013 13506 13030 13523
rect 14531 13506 14548 13523
rect 26215 13506 26232 13523
rect 3326 13472 3343 13489
rect 3481 13472 3498 13489
rect 4614 13472 4631 13489
rect 4706 13472 4723 13489
rect 4816 13472 4833 13489
rect 5166 13472 5183 13489
rect 5212 13472 5229 13489
rect 9168 13472 9185 13489
rect 9260 13472 9277 13489
rect 10203 13472 10220 13489
rect 12342 13472 12359 13489
rect 12434 13472 12451 13489
rect 12957 13472 12974 13489
rect 14475 13472 14492 13489
rect 15742 13472 15759 13489
rect 18414 13472 18431 13489
rect 18461 13472 18478 13489
rect 18832 13472 18849 13489
rect 19058 13472 19075 13489
rect 24210 13472 24227 13489
rect 26004 13472 26021 13489
rect 26159 13472 26176 13489
rect 4752 13438 4769 13455
rect 6914 13438 6931 13455
rect 10042 13438 10059 13455
rect 12802 13438 12819 13455
rect 14320 13438 14337 13455
rect 15608 13438 15625 13455
rect 18966 13438 18983 13455
rect 24164 13438 24181 13455
rect 24302 13438 24319 13455
rect 9214 13404 9231 13421
rect 9490 13404 9507 13421
rect 18598 13404 18615 13421
rect 19012 13404 19029 13421
rect 5212 13370 5229 13387
rect 7949 13370 7966 13387
rect 9766 13370 9783 13387
rect 11077 13370 11094 13387
rect 12388 13370 12405 13387
rect 13837 13370 13854 13387
rect 18897 13370 18914 13387
rect 24256 13370 24273 13387
rect 4177 13268 4194 13285
rect 12457 13268 12474 13285
rect 16068 13268 16085 13285
rect 18782 13268 18799 13285
rect 7880 13234 7897 13251
rect 16344 13234 16361 13251
rect 3142 13200 3159 13217
rect 4798 13200 4815 13217
rect 5350 13200 5367 13217
rect 11422 13200 11439 13217
rect 15976 13200 15993 13217
rect 16114 13200 16131 13217
rect 3303 13166 3320 13183
rect 4752 13166 4769 13183
rect 4847 13166 4864 13183
rect 7880 13166 7897 13183
rect 7937 13166 7954 13183
rect 8031 13164 8048 13181
rect 8093 13166 8110 13183
rect 8141 13156 8158 13173
rect 8192 13166 8209 13183
rect 8662 13166 8679 13183
rect 11577 13166 11594 13183
rect 13262 13166 13279 13183
rect 14550 13166 14567 13183
rect 14627 13166 14644 13183
rect 14701 13164 14718 13181
rect 14749 13172 14766 13189
rect 14811 13172 14828 13189
rect 14862 13166 14879 13183
rect 16022 13166 16039 13183
rect 16344 13166 16361 13183
rect 16482 13166 16499 13183
rect 18644 13166 18661 13183
rect 18736 13166 18753 13183
rect 18782 13166 18799 13183
rect 21220 13166 21237 13183
rect 21381 13166 21398 13183
rect 3353 13132 3370 13149
rect 4660 13132 4677 13149
rect 4798 13132 4815 13149
rect 5511 13132 5528 13149
rect 5561 13132 5578 13149
rect 8822 13132 8839 13149
rect 8873 13132 8890 13149
rect 11633 13132 11650 13149
rect 13422 13132 13439 13149
rect 13473 13132 13490 13149
rect 21431 13132 21448 13149
rect 6385 13098 6402 13115
rect 9697 13098 9714 13115
rect 14297 13098 14314 13115
rect 14550 13098 14567 13115
rect 16436 13098 16453 13115
rect 22255 13098 22272 13115
rect 4683 12996 4700 13013
rect 7995 12996 8012 13013
rect 11974 12996 11991 13013
rect 12342 12996 12359 13013
rect 12388 12996 12405 13013
rect 13837 12996 13854 13013
rect 19334 12996 19351 13013
rect 29500 12996 29517 13013
rect 3859 12962 3876 12979
rect 6316 12962 6333 12979
rect 6362 12962 6379 12979
rect 7171 12962 7188 12979
rect 10249 12962 10266 12979
rect 11077 12962 11094 12979
rect 13013 12962 13030 12979
rect 19242 12962 19259 12979
rect 20966 12962 20983 12979
rect 21017 12962 21034 12979
rect 26073 12962 26090 12979
rect 28372 12962 28389 12979
rect 28423 12962 28440 12979
rect 3809 12928 3826 12945
rect 6178 12928 6195 12945
rect 6224 12928 6241 12945
rect 6408 12928 6425 12945
rect 7115 12928 7132 12945
rect 10203 12928 10220 12945
rect 11744 12928 11761 12945
rect 11801 12928 11818 12945
rect 11895 12928 11912 12945
rect 11957 12923 11974 12940
rect 12005 12923 12022 12940
rect 12056 12928 12073 12945
rect 12296 12928 12313 12945
rect 12480 12928 12497 12945
rect 12957 12928 12974 12945
rect 16160 12928 16177 12945
rect 16482 12928 16499 12945
rect 19196 12928 19213 12945
rect 19380 12928 19397 12945
rect 21841 12928 21858 12945
rect 22600 12928 22617 12945
rect 22657 12928 22674 12945
rect 22751 12931 22768 12948
rect 22813 12923 22830 12940
rect 22861 12923 22878 12940
rect 22912 12928 22929 12945
rect 26027 12928 26044 12945
rect 29500 12928 29517 12945
rect 29557 12928 29574 12945
rect 29661 12928 29678 12945
rect 29713 12928 29730 12945
rect 29761 12928 29778 12945
rect 29812 12928 29829 12945
rect 3648 12894 3665 12911
rect 6454 12894 6471 12911
rect 6960 12894 6977 12911
rect 10042 12894 10059 12911
rect 12802 12894 12819 12911
rect 16528 12894 16545 12911
rect 19288 12894 19305 12911
rect 20806 12894 20823 12911
rect 25866 12894 25883 12911
rect 28212 12894 28229 12911
rect 29247 12894 29264 12911
rect 12434 12826 12451 12843
rect 22600 12826 22617 12843
rect 26901 12826 26918 12843
rect 4177 12724 4194 12741
rect 6247 12724 6264 12741
rect 9145 12724 9162 12741
rect 11905 12724 11922 12741
rect 13998 12724 14015 12741
rect 22255 12724 22272 12741
rect 28879 12724 28896 12741
rect 3142 12656 3159 12673
rect 5212 12656 5229 12673
rect 8110 12656 8127 12673
rect 10870 12656 10887 12673
rect 21220 12656 21237 12673
rect 3303 12622 3320 12639
rect 5411 12622 5428 12639
rect 6500 12622 6517 12639
rect 6638 12622 6655 12639
rect 11025 12622 11042 12639
rect 14504 12622 14521 12639
rect 14550 12622 14567 12639
rect 14688 12622 14705 12639
rect 15700 12622 15717 12639
rect 15792 12622 15809 12639
rect 16436 12622 16453 12639
rect 16528 12622 16545 12639
rect 16758 12622 16775 12639
rect 20070 12622 20087 12639
rect 20300 12622 20317 12639
rect 21375 12622 21392 12639
rect 21419 12622 21436 12639
rect 27844 12622 27861 12639
rect 28005 12622 28022 12639
rect 3353 12588 3370 12605
rect 5372 12588 5389 12605
rect 6592 12588 6609 12605
rect 8270 12588 8287 12605
rect 8321 12588 8338 12605
rect 11081 12588 11098 12605
rect 13906 12588 13923 12605
rect 20438 12588 20455 12605
rect 28055 12588 28072 12605
rect 6546 12554 6563 12571
rect 14006 12554 14023 12571
rect 14090 12554 14107 12571
rect 14596 12554 14613 12571
rect 14688 12554 14705 12571
rect 15746 12554 15763 12571
rect 12120 12452 12137 12469
rect 12204 12452 12221 12469
rect 23980 12452 23997 12469
rect 27154 12452 27171 12469
rect 4733 12418 4750 12435
rect 7075 12418 7092 12435
rect 8960 12418 8977 12435
rect 9011 12418 9028 12435
rect 12020 12418 12037 12435
rect 12779 12418 12796 12435
rect 14480 12418 14497 12435
rect 14531 12418 14548 12435
rect 15742 12418 15759 12435
rect 17080 12418 17097 12435
rect 18322 12418 18339 12435
rect 18414 12418 18431 12435
rect 25571 12418 25588 12435
rect 27338 12418 27355 12435
rect 28280 12418 28297 12435
rect 28331 12418 28348 12435
rect 4683 12384 4700 12401
rect 6868 12384 6885 12401
rect 7029 12384 7046 12401
rect 7903 12384 7920 12401
rect 8800 12384 8817 12401
rect 10088 12384 10105 12401
rect 11560 12384 11577 12401
rect 11652 12384 11669 12401
rect 11698 12384 11715 12401
rect 11747 12384 11764 12401
rect 12733 12384 12750 12401
rect 15608 12384 15625 12401
rect 17172 12384 17189 12401
rect 17218 12384 17235 12401
rect 17267 12379 17284 12396
rect 17770 12384 17787 12401
rect 17862 12384 17879 12401
rect 17908 12384 17925 12401
rect 18460 12384 18477 12401
rect 19150 12384 19167 12401
rect 19242 12384 19259 12401
rect 19288 12384 19305 12401
rect 23888 12384 23905 12401
rect 23934 12384 23951 12401
rect 25360 12384 25377 12401
rect 25521 12384 25538 12401
rect 26395 12384 26412 12401
rect 26648 12384 26665 12401
rect 26740 12384 26757 12401
rect 26786 12384 26803 12401
rect 26832 12384 26849 12401
rect 27154 12384 27171 12401
rect 27200 12384 27217 12401
rect 27292 12384 27309 12401
rect 27384 12384 27401 12401
rect 29155 12384 29172 12401
rect 4522 12350 4539 12367
rect 10870 12350 10887 12367
rect 11606 12350 11623 12367
rect 12572 12350 12589 12367
rect 14320 12350 14337 12367
rect 24072 12350 24089 12367
rect 28120 12350 28137 12367
rect 19288 12316 19305 12333
rect 26924 12316 26941 12333
rect 5557 12282 5574 12299
rect 9835 12282 9852 12299
rect 12112 12282 12129 12299
rect 13607 12282 13624 12299
rect 15355 12282 15372 12299
rect 16298 12282 16315 12299
rect 17080 12282 17097 12299
rect 17816 12282 17833 12299
rect 18460 12282 18477 12299
rect 23934 12282 23951 12299
rect 7420 12180 7437 12197
rect 11215 12180 11232 12197
rect 14228 12180 14245 12197
rect 14872 12180 14889 12197
rect 15792 12180 15809 12197
rect 16988 12180 17005 12197
rect 19932 12180 19949 12197
rect 26257 12180 26274 12197
rect 5580 12146 5597 12163
rect 19518 12146 19535 12163
rect 22002 12146 22019 12163
rect 4706 12112 4723 12129
rect 6845 12112 6862 12129
rect 8528 12112 8545 12129
rect 10180 12112 10197 12129
rect 11974 12112 11991 12129
rect 16229 12112 16246 12129
rect 18506 12112 18523 12129
rect 18736 12112 18753 12129
rect 19840 12112 19857 12129
rect 19978 12112 19995 12129
rect 25222 12112 25239 12129
rect 5810 12078 5827 12095
rect 5965 12078 5982 12095
rect 7420 12078 7437 12095
rect 7466 12078 7483 12095
rect 7558 12078 7575 12095
rect 7604 12078 7621 12095
rect 7650 12078 7667 12095
rect 10341 12078 10358 12095
rect 12023 12078 12040 12095
rect 12940 12078 12957 12095
rect 14228 12078 14245 12095
rect 14320 12078 14337 12095
rect 14415 12078 14432 12095
rect 14826 12078 14843 12095
rect 14918 12078 14935 12095
rect 15930 12078 15947 12095
rect 16178 12078 16195 12095
rect 16988 12078 17005 12095
rect 17080 12078 17097 12095
rect 17402 12078 17419 12095
rect 17540 12078 17557 12095
rect 18552 12078 18569 12095
rect 19472 12078 19489 12095
rect 19886 12078 19903 12095
rect 21956 12078 21973 12095
rect 22094 12078 22111 12095
rect 25383 12078 25400 12095
rect 4844 12044 4861 12061
rect 6021 12044 6038 12061
rect 8684 12044 8701 12061
rect 8735 12044 8752 12061
rect 10391 12044 10408 12061
rect 11836 12044 11853 12061
rect 11928 12044 11945 12061
rect 11974 12044 11991 12061
rect 13100 12044 13117 12061
rect 13151 12044 13168 12061
rect 14366 12044 14383 12061
rect 15792 12044 15809 12061
rect 15884 12044 15901 12061
rect 19610 12044 19627 12061
rect 22048 12044 22065 12061
rect 25433 12044 25450 12061
rect 9559 12010 9576 12027
rect 13975 12010 13992 12027
rect 17448 12010 17465 12027
rect 19472 12010 19489 12027
rect 5212 11908 5229 11925
rect 5396 11908 5413 11925
rect 5442 11908 5459 11925
rect 9214 11908 9231 11925
rect 10985 11908 11002 11925
rect 16114 11908 16131 11925
rect 19380 11908 19397 11925
rect 26947 11908 26964 11925
rect 7489 11874 7506 11891
rect 8317 11874 8334 11891
rect 9076 11874 9093 11891
rect 9628 11874 9645 11891
rect 10157 11874 10174 11891
rect 13013 11874 13030 11891
rect 13837 11874 13854 11891
rect 14458 11874 14475 11891
rect 20419 11874 20436 11891
rect 26072 11874 26089 11891
rect 26123 11874 26140 11891
rect 6086 11840 6103 11857
rect 7443 11840 7460 11857
rect 8938 11840 8955 11857
rect 9030 11840 9047 11857
rect 9122 11840 9139 11857
rect 9444 11840 9461 11857
rect 9490 11840 9507 11857
rect 9582 11840 9599 11857
rect 9674 11840 9691 11857
rect 10111 11840 10128 11857
rect 11882 11840 11899 11857
rect 12802 11840 12819 11857
rect 12957 11840 12974 11857
rect 14320 11840 14337 11857
rect 14412 11840 14429 11857
rect 14507 11840 14524 11857
rect 16114 11840 16131 11857
rect 16252 11840 16269 11857
rect 16298 11840 16315 11857
rect 18690 11840 18707 11857
rect 18818 11840 18835 11857
rect 20363 11840 20380 11857
rect 21243 11840 21260 11857
rect 21542 11840 21559 11857
rect 21634 11840 21651 11857
rect 21680 11840 21697 11857
rect 21729 11840 21746 11857
rect 25912 11840 25929 11857
rect 5488 11806 5505 11823
rect 6868 11806 6885 11823
rect 7052 11806 7069 11823
rect 7282 11806 7299 11823
rect 9720 11806 9737 11823
rect 9950 11806 9967 11823
rect 12388 11806 12405 11823
rect 20208 11806 20225 11823
rect 21588 11806 21605 11823
rect 14320 11772 14337 11789
rect 7696 11636 7713 11653
rect 9697 11636 9714 11653
rect 11997 11636 12014 11653
rect 13975 11636 13992 11653
rect 18690 11636 18707 11653
rect 8662 11568 8679 11585
rect 12940 11568 12957 11585
rect 16482 11568 16499 11585
rect 5902 11534 5919 11551
rect 6063 11534 6080 11551
rect 6937 11534 6954 11551
rect 7420 11534 7437 11551
rect 7512 11534 7529 11551
rect 7604 11534 7621 11551
rect 8861 11534 8878 11551
rect 10272 11534 10289 11551
rect 10318 11534 10335 11551
rect 10962 11534 10979 11551
rect 11117 11534 11134 11551
rect 16344 11534 16361 11551
rect 16390 11534 16407 11551
rect 18644 11534 18661 11551
rect 18736 11534 18753 11551
rect 19472 11534 19489 11551
rect 19564 11534 19581 11551
rect 6113 11500 6130 11517
rect 7558 11500 7575 11517
rect 8822 11500 8839 11517
rect 10180 11500 10197 11517
rect 11173 11500 11190 11517
rect 13100 11500 13117 11517
rect 13151 11500 13168 11517
rect 19610 11500 19627 11517
rect 10318 11466 10335 11483
rect 16344 11466 16361 11483
rect 21519 11364 21536 11381
rect 24440 11364 24457 11381
rect 4733 11330 4750 11347
rect 6752 11330 6769 11347
rect 6803 11330 6820 11347
rect 17494 11330 17511 11347
rect 20695 11330 20712 11347
rect 28331 11330 28348 11347
rect 29155 11330 29172 11347
rect 4522 11296 4539 11313
rect 4683 11296 4700 11313
rect 16206 11296 16223 11313
rect 16298 11296 16315 11313
rect 17126 11296 17143 11313
rect 17448 11296 17465 11313
rect 17540 11296 17557 11313
rect 18460 11296 18477 11313
rect 18552 11296 18569 11313
rect 20639 11296 20656 11313
rect 24348 11296 24365 11313
rect 24486 11296 24503 11313
rect 24578 11296 24595 11313
rect 28281 11296 28298 11313
rect 29408 11296 29425 11313
rect 29500 11296 29517 11313
rect 6592 11262 6609 11279
rect 7627 11262 7644 11279
rect 17080 11262 17097 11279
rect 17218 11262 17235 11279
rect 20484 11262 20501 11279
rect 28120 11262 28137 11279
rect 16068 11228 16085 11245
rect 17172 11228 17189 11245
rect 5557 11194 5574 11211
rect 16206 11194 16223 11211
rect 18506 11194 18523 11211
rect 29454 11194 29471 11211
rect 18460 11092 18477 11109
rect 6661 11058 6678 11075
rect 16942 11058 16959 11075
rect 5350 11024 5367 11041
rect 11859 11024 11876 11041
rect 13952 11024 13969 11041
rect 16344 11024 16361 11041
rect 17218 11024 17235 11041
rect 21220 11024 21237 11041
rect 22508 11024 22525 11041
rect 5258 10990 5275 11007
rect 5626 10990 5643 11007
rect 5781 10990 5798 11007
rect 10824 10990 10841 11007
rect 10985 10990 11002 11007
rect 16206 10990 16223 11007
rect 16252 10990 16269 11007
rect 16390 10990 16407 11007
rect 16896 10990 16913 11007
rect 17172 10990 17189 11007
rect 18460 10990 18477 11007
rect 18598 10990 18615 11007
rect 22695 10990 22712 11007
rect 23152 10990 23169 11007
rect 23244 10990 23261 11007
rect 23980 10990 23997 11007
rect 24072 10990 24089 11007
rect 5837 10956 5854 10973
rect 11035 10956 11052 10973
rect 18552 10956 18569 10973
rect 21380 10956 21397 10973
rect 21431 10956 21448 10973
rect 22255 10956 22272 10973
rect 22508 10956 22525 10973
rect 22600 10956 22617 10973
rect 22646 10956 22663 10973
rect 5028 10922 5045 10939
rect 5212 10922 5229 10939
rect 13676 10922 13693 10939
rect 13860 10922 13877 10939
rect 13906 10922 13923 10939
rect 16114 10922 16131 10939
rect 23198 10922 23215 10939
rect 24026 10922 24043 10939
rect 13423 10820 13440 10837
rect 15792 10820 15809 10837
rect 22117 10820 22134 10837
rect 22968 10820 22985 10837
rect 26832 10820 26849 10837
rect 29086 10820 29103 10837
rect 10249 10786 10266 10803
rect 11077 10786 11094 10803
rect 12548 10786 12565 10803
rect 12599 10786 12616 10803
rect 14669 10786 14686 10803
rect 15493 10786 15510 10803
rect 20208 10786 20225 10803
rect 21281 10786 21298 10803
rect 23367 10786 23384 10803
rect 24287 10786 24304 10803
rect 25571 10786 25588 10803
rect 29132 10786 29149 10803
rect 10042 10752 10059 10769
rect 10203 10752 10220 10769
rect 11836 10752 11853 10769
rect 12158 10752 12175 10769
rect 14619 10752 14636 10769
rect 15792 10752 15809 10769
rect 16206 10752 16223 10769
rect 18276 10752 18293 10769
rect 18818 10752 18835 10769
rect 20300 10752 20317 10769
rect 20346 10752 20363 10769
rect 21237 10752 21254 10769
rect 22922 10752 22939 10769
rect 23014 10752 23031 10769
rect 25521 10752 25538 10769
rect 26694 10752 26711 10769
rect 29040 10752 29057 10769
rect 29178 10752 29195 10769
rect 11928 10718 11945 10735
rect 12388 10718 12405 10735
rect 14458 10718 14475 10735
rect 18322 10718 18339 10735
rect 18690 10718 18707 10735
rect 21082 10718 21099 10735
rect 23244 10718 23261 10735
rect 24164 10718 24181 10735
rect 25360 10718 25377 10735
rect 26832 10718 26849 10735
rect 19380 10684 19397 10701
rect 18414 10650 18431 10667
rect 20208 10650 20225 10667
rect 23934 10650 23951 10667
rect 24854 10650 24871 10667
rect 26395 10650 26412 10667
rect 26740 10650 26757 10667
rect 17172 10548 17189 10565
rect 18690 10548 18707 10565
rect 20415 10548 20432 10565
rect 23014 10548 23031 10565
rect 23428 10548 23445 10565
rect 24072 10548 24089 10565
rect 14780 10514 14797 10531
rect 4982 10480 4999 10497
rect 5120 10480 5137 10497
rect 8432 10480 8449 10497
rect 8754 10480 8771 10497
rect 13676 10480 13693 10497
rect 14550 10480 14567 10497
rect 16022 10480 16039 10497
rect 19380 10480 19397 10497
rect 23474 10480 23491 10497
rect 24118 10480 24135 10497
rect 24624 10480 24641 10497
rect 25659 10480 25676 10497
rect 28948 10480 28965 10497
rect 8340 10446 8357 10463
rect 8524 10446 8541 10463
rect 13538 10446 13555 10463
rect 14918 10446 14935 10463
rect 15884 10446 15901 10463
rect 17218 10446 17235 10463
rect 17402 10446 17419 10463
rect 18644 10446 18661 10463
rect 18736 10446 18753 10463
rect 19541 10446 19558 10463
rect 23014 10446 23031 10463
rect 23106 10446 23123 10463
rect 23336 10446 23353 10463
rect 23382 10446 23399 10463
rect 23980 10446 23997 10463
rect 24026 10446 24043 10463
rect 24785 10446 24802 10463
rect 25912 10446 25929 10463
rect 25969 10446 25986 10463
rect 26063 10446 26080 10463
rect 26111 10452 26128 10469
rect 26173 10444 26190 10461
rect 26224 10446 26241 10463
rect 27522 10446 27539 10463
rect 28902 10446 28919 10463
rect 28997 10446 29014 10463
rect 5994 10412 6011 10429
rect 8892 10412 8909 10429
rect 14780 10412 14797 10429
rect 16896 10412 16913 10429
rect 19591 10412 19608 10429
rect 24831 10412 24848 10429
rect 27682 10412 27699 10429
rect 27733 10412 27750 10429
rect 28557 10412 28574 10429
rect 28810 10412 28827 10429
rect 28948 10412 28965 10429
rect 8386 10378 8403 10395
rect 8478 10378 8495 10395
rect 9628 10378 9645 10395
rect 14872 10378 14889 10395
rect 26142 10378 26159 10395
rect 26395 10276 26412 10293
rect 29155 10276 29172 10293
rect 9030 10242 9047 10259
rect 14454 10242 14471 10259
rect 15746 10242 15763 10259
rect 25571 10242 25588 10259
rect 28331 10242 28348 10259
rect 8064 10208 8081 10225
rect 8846 10208 8863 10225
rect 8938 10208 8955 10225
rect 9536 10208 9553 10225
rect 15608 10208 15625 10225
rect 25360 10208 25377 10225
rect 25521 10208 25538 10225
rect 28120 10208 28137 10225
rect 28281 10208 28298 10225
rect 8018 10174 8035 10191
rect 9674 10174 9691 10191
rect 10548 10174 10565 10191
rect 14320 10174 14337 10191
rect 16620 10174 16637 10191
rect 8202 10106 8219 10123
rect 15010 10106 15027 10123
rect 7512 10004 7529 10021
rect 9122 10004 9139 10021
rect 9674 10004 9691 10021
rect 19150 9970 19167 9987
rect 7926 9936 7943 9953
rect 8800 9936 8817 9953
rect 9214 9936 9231 9953
rect 9582 9936 9599 9953
rect 10180 9936 10197 9953
rect 14366 9936 14383 9953
rect 14504 9936 14521 9953
rect 17494 9936 17511 9953
rect 17908 9936 17925 9953
rect 18000 9936 18017 9953
rect 22278 9936 22295 9953
rect 7466 9902 7483 9919
rect 7558 9902 7575 9919
rect 7788 9902 7805 9919
rect 9168 9902 9185 9919
rect 9536 9902 9553 9919
rect 14412 9902 14429 9919
rect 17126 9902 17143 9919
rect 17356 9902 17373 9919
rect 17862 9902 17879 9919
rect 18460 9902 18477 9919
rect 22508 9902 22525 9919
rect 9030 9868 9047 9885
rect 10318 9868 10335 9885
rect 14504 9868 14521 9885
rect 18583 9868 18600 9885
rect 22324 9868 22341 9885
rect 22554 9868 22571 9885
rect 22600 9868 22617 9885
rect 9076 9834 9093 9851
rect 11054 9834 11071 9851
rect 17172 9834 17189 9851
rect 17862 9834 17879 9851
rect 8892 9732 8909 9749
rect 8984 9732 9001 9749
rect 14458 9732 14475 9749
rect 20622 9732 20639 9749
rect 23428 9732 23445 9749
rect 8846 9698 8863 9715
rect 9490 9698 9507 9715
rect 14366 9698 14383 9715
rect 17172 9698 17189 9715
rect 19196 9698 19213 9715
rect 7926 9664 7943 9681
rect 8800 9664 8817 9681
rect 9582 9664 9599 9681
rect 9996 9664 10013 9681
rect 14504 9664 14521 9681
rect 17080 9664 17097 9681
rect 19104 9664 19121 9681
rect 19150 9664 19167 9681
rect 20530 9664 20547 9681
rect 20576 9664 20593 9681
rect 22600 9664 22617 9681
rect 22692 9664 22709 9681
rect 23106 9664 23123 9681
rect 23336 9664 23353 9681
rect 7880 9630 7897 9647
rect 8984 9630 9001 9647
rect 9674 9630 9691 9647
rect 9950 9630 9967 9647
rect 10180 9630 10197 9647
rect 17264 9630 17281 9647
rect 19012 9630 19029 9647
rect 19380 9630 19397 9647
rect 20714 9630 20731 9647
rect 8846 9596 8863 9613
rect 20576 9596 20593 9613
rect 8110 9562 8127 9579
rect 14366 9562 14383 9579
rect 15056 9460 15073 9477
rect 20530 9460 20547 9477
rect 27016 9460 27033 9477
rect 29500 9460 29517 9477
rect 7788 9392 7805 9409
rect 8662 9392 8679 9409
rect 15010 9392 15027 9409
rect 15102 9392 15119 9409
rect 23980 9392 23997 9409
rect 25268 9392 25285 9409
rect 27154 9392 27171 9409
rect 27982 9392 27999 9409
rect 7650 9358 7667 9375
rect 14044 9358 14061 9375
rect 14178 9358 14195 9375
rect 14964 9358 14981 9375
rect 15884 9358 15901 9375
rect 18874 9358 18891 9375
rect 18966 9358 18983 9375
rect 19380 9358 19397 9375
rect 19610 9358 19627 9375
rect 20622 9358 20639 9375
rect 20668 9358 20685 9375
rect 20732 9358 20749 9375
rect 22140 9358 22157 9375
rect 22232 9358 22249 9375
rect 22646 9358 22663 9375
rect 22876 9358 22893 9375
rect 25455 9358 25472 9375
rect 26970 9358 26987 9375
rect 29592 9358 29609 9375
rect 29687 9358 29704 9375
rect 15746 9324 15763 9341
rect 15838 9324 15855 9341
rect 20530 9324 20547 9341
rect 24140 9324 24157 9341
rect 24191 9324 24208 9341
rect 25015 9324 25032 9341
rect 25268 9324 25285 9341
rect 25360 9324 25377 9341
rect 25406 9324 25423 9341
rect 28142 9324 28159 9341
rect 28193 9324 28210 9341
rect 29017 9324 29034 9341
rect 29500 9324 29517 9341
rect 29638 9324 29655 9341
rect 14734 9290 14751 9307
rect 15792 9290 15809 9307
rect 19058 9290 19075 9307
rect 19702 9290 19719 9307
rect 22968 9290 22985 9307
rect 27016 9290 27033 9307
rect 27062 9290 27079 9307
rect 14734 9188 14751 9205
rect 20875 9188 20892 9205
rect 22784 9188 22801 9205
rect 23428 9188 23445 9205
rect 24877 9188 24894 9205
rect 26924 9188 26941 9205
rect 29155 9188 29172 9205
rect 19288 9154 19305 9171
rect 20051 9154 20068 9171
rect 24041 9154 24058 9171
rect 25796 9154 25813 9171
rect 25847 9154 25864 9171
rect 28280 9154 28297 9171
rect 28331 9154 28348 9171
rect 13768 9120 13785 9137
rect 13860 9120 13877 9137
rect 14550 9120 14567 9137
rect 15286 9120 15303 9137
rect 16058 9120 16075 9137
rect 18966 9120 18983 9137
rect 19196 9120 19213 9137
rect 19242 9120 19259 9137
rect 20001 9120 20018 9137
rect 22600 9120 22617 9137
rect 22692 9120 22709 9137
rect 23106 9120 23123 9137
rect 23336 9120 23353 9137
rect 23997 9120 24014 9137
rect 26924 9120 26941 9137
rect 26981 9120 26998 9137
rect 27082 9120 27099 9137
rect 27130 9120 27147 9137
rect 27185 9120 27202 9137
rect 27236 9120 27253 9137
rect 28120 9120 28137 9137
rect 14596 9086 14613 9103
rect 15240 9086 15257 9103
rect 15470 9086 15487 9103
rect 15930 9086 15947 9103
rect 17080 9086 17097 9103
rect 17126 9086 17143 9103
rect 17218 9086 17235 9103
rect 19012 9086 19029 9103
rect 19840 9086 19857 9103
rect 23842 9086 23859 9103
rect 25636 9086 25653 9103
rect 26671 9086 26688 9103
rect 14734 9052 14751 9069
rect 16620 9052 16637 9069
rect 13768 9018 13785 9035
rect 17172 9018 17189 9035
rect 14504 8916 14521 8933
rect 15976 8916 15993 8933
rect 17862 8916 17879 8933
rect 20737 8916 20754 8933
rect 27775 8916 27792 8933
rect 7788 8882 7805 8899
rect 14136 8882 14153 8899
rect 5902 8848 5919 8865
rect 6040 8848 6057 8865
rect 7696 8848 7713 8865
rect 10364 8848 10381 8865
rect 11376 8848 11393 8865
rect 14596 8848 14613 8865
rect 19702 8848 19719 8865
rect 26740 8848 26757 8865
rect 5856 8814 5873 8831
rect 7604 8814 7621 8831
rect 7788 8814 7805 8831
rect 8018 8814 8035 8831
rect 8110 8814 8127 8831
rect 13446 8814 13463 8831
rect 13580 8814 13597 8831
rect 14412 8814 14429 8831
rect 14550 8814 14567 8831
rect 15792 8814 15809 8831
rect 15838 8814 15855 8831
rect 15884 8814 15901 8831
rect 18000 8814 18017 8831
rect 19863 8814 19880 8831
rect 22186 8814 22203 8831
rect 22278 8814 22295 8831
rect 22554 8814 22571 8831
rect 22830 8814 22847 8831
rect 10502 8780 10519 8797
rect 14366 8780 14383 8797
rect 15700 8780 15717 8797
rect 15976 8780 15993 8797
rect 17862 8780 17879 8797
rect 19913 8780 19930 8797
rect 26901 8780 26918 8797
rect 26951 8780 26968 8797
rect 7650 8746 7667 8763
rect 8064 8746 8081 8763
rect 17954 8746 17971 8763
rect 22738 8746 22755 8763
rect 7742 8644 7759 8661
rect 9536 8644 9553 8661
rect 10502 8644 10519 8661
rect 18414 8644 18431 8661
rect 22876 8644 22893 8661
rect 26855 8644 26872 8661
rect 7834 8610 7851 8627
rect 8018 8610 8035 8627
rect 9214 8610 9231 8627
rect 10686 8610 10703 8627
rect 23589 8610 23606 8627
rect 26027 8610 26044 8627
rect 28810 8610 28827 8627
rect 28856 8610 28873 8627
rect 7788 8576 7805 8593
rect 9076 8576 9093 8593
rect 9490 8576 9507 8593
rect 10456 8576 10473 8593
rect 10916 8576 10933 8593
rect 11008 8576 11025 8593
rect 17080 8576 17097 8593
rect 17172 8576 17189 8593
rect 18230 8576 18247 8593
rect 21266 8576 21283 8593
rect 21450 8576 21467 8593
rect 21634 8576 21651 8593
rect 22048 8576 22065 8593
rect 22600 8576 22617 8593
rect 22738 8576 22755 8593
rect 22876 8576 22893 8593
rect 23382 8576 23399 8593
rect 23537 8576 23554 8593
rect 25975 8576 25992 8593
rect 28718 8576 28735 8593
rect 28905 8576 28922 8593
rect 6408 8542 6425 8559
rect 6546 8542 6563 8559
rect 7420 8542 7437 8559
rect 7650 8542 7667 8559
rect 8938 8542 8955 8559
rect 9168 8542 9185 8559
rect 10640 8542 10657 8559
rect 18276 8542 18293 8559
rect 22968 8542 22985 8559
rect 25820 8542 25837 8559
rect 9030 8508 9047 8525
rect 10594 8508 10611 8525
rect 10916 8508 10933 8525
rect 17218 8508 17235 8525
rect 21818 8508 21835 8525
rect 23106 8508 23123 8525
rect 28718 8508 28735 8525
rect 8984 8474 9001 8491
rect 24417 8474 24434 8491
rect 8524 8372 8541 8389
rect 8938 8372 8955 8389
rect 5856 8304 5873 8321
rect 7788 8304 7805 8321
rect 5718 8270 5735 8287
rect 6730 8270 6747 8287
rect 7650 8270 7667 8287
rect 9398 8270 9415 8287
rect 19610 8270 19627 8287
rect 19794 8270 19811 8287
rect 19840 8270 19857 8287
rect 19932 8270 19949 8287
rect 22140 8270 22157 8287
rect 22232 8270 22249 8287
rect 22738 8270 22755 8287
rect 22876 8270 22893 8287
rect 24256 8270 24273 8287
rect 24333 8270 24350 8287
rect 24407 8268 24424 8285
rect 24469 8270 24486 8287
rect 24517 8268 24534 8285
rect 24568 8268 24585 8285
rect 8800 8236 8817 8253
rect 8846 8202 8863 8219
rect 22968 8202 22985 8219
rect 24486 8202 24503 8219
rect 15516 8100 15533 8117
rect 17356 8100 17373 8117
rect 18598 8100 18615 8117
rect 21358 8100 21375 8117
rect 24233 8100 24250 8117
rect 24762 8100 24779 8117
rect 24808 8100 24825 8117
rect 29155 8100 29172 8117
rect 20162 8066 20179 8083
rect 20392 8066 20409 8083
rect 20438 8066 20455 8083
rect 23409 8066 23426 8083
rect 28331 8066 28348 8083
rect 6408 8032 6425 8049
rect 6546 8032 6563 8049
rect 6638 8032 6655 8049
rect 8110 8032 8127 8049
rect 8202 8032 8219 8049
rect 8248 8032 8265 8049
rect 10732 8032 10749 8049
rect 14412 8032 14429 8049
rect 14504 8032 14521 8049
rect 14550 8032 14567 8049
rect 15332 8032 15349 8049
rect 17172 8032 17189 8049
rect 18414 8032 18431 8049
rect 20116 8032 20133 8049
rect 20346 8032 20363 8049
rect 20806 8032 20823 8049
rect 21082 8032 21099 8049
rect 21174 8032 21191 8049
rect 21542 8032 21559 8049
rect 23198 8032 23215 8049
rect 23359 8032 23376 8049
rect 24716 8032 24733 8049
rect 24900 8032 24917 8049
rect 28281 8032 28298 8049
rect 6868 7998 6885 8015
rect 7006 7998 7023 8015
rect 7880 7998 7897 8015
rect 10870 7998 10887 8015
rect 15286 7998 15303 8015
rect 17126 7998 17143 8015
rect 17402 7998 17419 8015
rect 18460 7998 18477 8015
rect 28120 7998 28137 8015
rect 6408 7964 6425 7981
rect 10778 7964 10795 7981
rect 17356 7964 17373 7981
rect 24762 7964 24779 7981
rect 6546 7930 6563 7947
rect 8110 7930 8127 7947
rect 10732 7930 10749 7947
rect 14320 7930 14337 7947
rect 6822 7828 6839 7845
rect 7604 7828 7621 7845
rect 15976 7828 15993 7845
rect 17494 7828 17511 7845
rect 28971 7828 28988 7845
rect 29500 7828 29517 7845
rect 7650 7794 7667 7811
rect 26740 7794 26757 7811
rect 10548 7760 10565 7777
rect 10686 7760 10703 7777
rect 14136 7760 14153 7777
rect 15746 7760 15763 7777
rect 17402 7760 17419 7777
rect 19426 7760 19443 7777
rect 21542 7760 21559 7777
rect 6822 7726 6839 7743
rect 6960 7726 6977 7743
rect 7420 7726 7437 7743
rect 7650 7726 7667 7743
rect 13722 7726 13739 7743
rect 13814 7726 13831 7743
rect 13860 7726 13877 7743
rect 14090 7726 14107 7743
rect 14274 7726 14291 7743
rect 14366 7726 14383 7743
rect 15792 7726 15809 7743
rect 17356 7726 17373 7743
rect 19058 7726 19075 7743
rect 19288 7726 19305 7743
rect 19978 7726 19995 7743
rect 20116 7726 20133 7743
rect 21220 7726 21237 7743
rect 21450 7726 21467 7743
rect 22094 7726 22111 7743
rect 22186 7726 22203 7743
rect 22600 7726 22617 7743
rect 22830 7726 22847 7743
rect 26740 7726 26757 7743
rect 26817 7726 26834 7743
rect 26901 7716 26918 7733
rect 26953 7716 26970 7733
rect 27001 7726 27018 7743
rect 27052 7726 27069 7743
rect 27936 7726 27953 7743
rect 28091 7726 28108 7743
rect 29500 7726 29517 7743
rect 29546 7726 29563 7743
rect 29730 7726 29747 7743
rect 7466 7692 7483 7709
rect 11560 7692 11577 7709
rect 28135 7692 28152 7709
rect 29638 7692 29655 7709
rect 29684 7692 29701 7709
rect 6914 7658 6931 7675
rect 7512 7658 7529 7675
rect 8754 7658 8771 7675
rect 19932 7658 19949 7675
rect 22278 7658 22295 7675
rect 22922 7658 22939 7675
rect 6132 7556 6149 7573
rect 15516 7556 15533 7573
rect 18276 7556 18293 7573
rect 24325 7556 24342 7573
rect 26855 7556 26872 7573
rect 29155 7556 29172 7573
rect 6040 7522 6057 7539
rect 7144 7522 7161 7539
rect 8064 7522 8081 7539
rect 9352 7522 9369 7539
rect 9697 7522 9714 7539
rect 11652 7522 11669 7539
rect 19242 7522 19259 7539
rect 20484 7522 20501 7539
rect 20760 7522 20777 7539
rect 21036 7522 21053 7539
rect 21082 7522 21099 7539
rect 23497 7522 23514 7539
rect 26031 7522 26048 7539
rect 28331 7522 28348 7539
rect 6178 7488 6195 7505
rect 7926 7488 7943 7505
rect 9260 7488 9277 7505
rect 9398 7488 9415 7505
rect 9646 7488 9663 7505
rect 10410 7488 10427 7505
rect 10502 7488 10519 7505
rect 10732 7488 10749 7505
rect 10824 7488 10841 7505
rect 10870 7488 10887 7505
rect 11560 7488 11577 7505
rect 11698 7488 11715 7505
rect 15332 7488 15349 7505
rect 18230 7488 18247 7505
rect 18322 7488 18339 7505
rect 18966 7488 18983 7505
rect 19104 7488 19121 7505
rect 20116 7488 20133 7505
rect 20392 7488 20409 7505
rect 20990 7488 21007 7505
rect 23290 7488 23307 7505
rect 23451 7488 23468 7505
rect 25981 7488 25998 7505
rect 28120 7488 28137 7505
rect 28281 7488 28298 7505
rect 15286 7454 15303 7471
rect 20806 7454 20823 7471
rect 25820 7454 25837 7471
rect 7972 7420 7989 7437
rect 9260 7420 9277 7437
rect 11560 7420 11577 7437
rect 6040 7386 6057 7403
rect 7190 7386 7207 7403
rect 7926 7386 7943 7403
rect 10410 7386 10427 7403
rect 10732 7386 10749 7403
rect 10962 7386 10979 7403
rect 8846 7284 8863 7301
rect 9076 7284 9093 7301
rect 10769 7284 10786 7301
rect 14320 7284 14337 7301
rect 27775 7284 27792 7301
rect 12066 7250 12083 7267
rect 6546 7216 6563 7233
rect 7604 7216 7621 7233
rect 7742 7216 7759 7233
rect 8616 7216 8633 7233
rect 9720 7216 9737 7233
rect 10640 7216 10657 7233
rect 11652 7216 11669 7233
rect 12112 7216 12129 7233
rect 14090 7216 14107 7233
rect 19748 7216 19765 7233
rect 19840 7216 19857 7233
rect 26740 7216 26757 7233
rect 5534 7182 5551 7199
rect 8938 7182 8955 7199
rect 8984 7182 9001 7199
rect 9582 7182 9599 7199
rect 9628 7182 9645 7199
rect 11974 7182 11991 7199
rect 14136 7182 14153 7199
rect 18690 7182 18707 7199
rect 18828 7182 18845 7199
rect 18920 7182 18937 7199
rect 19564 7182 19581 7199
rect 19702 7182 19719 7199
rect 22232 7182 22249 7199
rect 22462 7182 22479 7199
rect 22646 7182 22663 7199
rect 22830 7182 22847 7199
rect 26895 7182 26912 7199
rect 5672 7148 5689 7165
rect 26951 7148 26968 7165
rect 9720 7114 9737 7131
rect 11882 7114 11899 7131
rect 18598 7114 18615 7131
rect 22370 7114 22387 7131
rect 6040 7012 6057 7029
rect 8294 7012 8311 7029
rect 11054 7012 11071 7029
rect 14458 7012 14475 7029
rect 20392 7012 20409 7029
rect 22117 7012 22134 7029
rect 10962 6978 10979 6995
rect 13722 6978 13739 6995
rect 13814 6978 13831 6995
rect 21293 6978 21310 6995
rect 23501 6978 23518 6995
rect 25893 6978 25910 6995
rect 29132 6978 29149 6995
rect 6132 6944 6149 6961
rect 8202 6944 8219 6961
rect 8340 6944 8357 6961
rect 11100 6944 11117 6961
rect 13860 6944 13877 6961
rect 14366 6944 14383 6961
rect 15792 6944 15809 6961
rect 16298 6944 16315 6961
rect 17954 6944 17971 6961
rect 18000 6944 18017 6961
rect 18092 6944 18109 6961
rect 18322 6944 18339 6961
rect 20116 6944 20133 6961
rect 20254 6944 20271 6961
rect 20346 6944 20363 6961
rect 21082 6944 21099 6961
rect 21237 6944 21254 6961
rect 22600 6944 22617 6961
rect 22657 6944 22674 6961
rect 22758 6944 22775 6961
rect 22806 6944 22823 6961
rect 22861 6955 22878 6972
rect 22912 6944 22929 6961
rect 23290 6944 23307 6961
rect 23451 6944 23468 6961
rect 24762 6944 24779 6961
rect 24854 6944 24871 6961
rect 24900 6944 24917 6961
rect 25843 6944 25860 6961
rect 29040 6944 29057 6961
rect 29178 6944 29195 6961
rect 29224 6944 29241 6961
rect 6270 6910 6287 6927
rect 14320 6910 14337 6927
rect 14458 6910 14475 6927
rect 15746 6910 15763 6927
rect 15976 6910 15993 6927
rect 16252 6910 16269 6927
rect 25682 6910 25699 6927
rect 8202 6876 8219 6893
rect 10962 6876 10979 6893
rect 16482 6876 16499 6893
rect 22600 6876 22617 6893
rect 24762 6876 24779 6893
rect 26717 6876 26734 6893
rect 29316 6876 29333 6893
rect 6224 6842 6241 6859
rect 13722 6842 13739 6859
rect 24325 6842 24342 6859
rect 14412 6740 14429 6757
rect 22255 6740 22272 6757
rect 25015 6740 25032 6757
rect 29017 6740 29034 6757
rect 6960 6672 6977 6689
rect 10824 6672 10841 6689
rect 10962 6672 10979 6689
rect 19288 6672 19305 6689
rect 23980 6672 23997 6689
rect 27982 6672 27999 6689
rect 6086 6638 6103 6655
rect 6822 6638 6839 6655
rect 6868 6638 6885 6655
rect 13722 6638 13739 6655
rect 13850 6638 13867 6655
rect 17862 6638 17879 6655
rect 17954 6638 17971 6655
rect 18966 6638 18983 6655
rect 19150 6638 19167 6655
rect 19564 6638 19581 6655
rect 19794 6638 19811 6655
rect 21220 6638 21237 6655
rect 21375 6638 21392 6655
rect 24135 6638 24152 6655
rect 28143 6638 28160 6655
rect 5948 6604 5965 6621
rect 11836 6604 11853 6621
rect 19932 6604 19949 6621
rect 21431 6604 21448 6621
rect 24191 6604 24208 6621
rect 28193 6604 28210 6621
rect 5997 6570 6014 6587
rect 6040 6570 6057 6587
rect 6822 6570 6839 6587
rect 17908 6570 17925 6587
rect 6132 6468 6149 6485
rect 22117 6468 22134 6485
rect 24716 6468 24733 6485
rect 6086 6434 6103 6451
rect 6730 6434 6747 6451
rect 16068 6434 16085 6451
rect 17264 6434 17281 6451
rect 19380 6434 19397 6451
rect 20576 6434 20593 6451
rect 21293 6434 21310 6451
rect 23363 6434 23380 6451
rect 24532 6434 24549 6451
rect 24578 6434 24595 6451
rect 28423 6434 28440 6451
rect 6040 6400 6057 6417
rect 6270 6400 6287 6417
rect 15976 6400 15993 6417
rect 16114 6400 16131 6417
rect 16528 6400 16545 6417
rect 16620 6400 16637 6417
rect 17126 6400 17143 6417
rect 17172 6400 17189 6417
rect 18138 6400 18155 6417
rect 18322 6400 18339 6417
rect 18414 6400 18431 6417
rect 19104 6400 19121 6417
rect 19242 6400 19259 6417
rect 20208 6400 20225 6417
rect 20438 6400 20455 6417
rect 21082 6400 21099 6417
rect 21243 6400 21260 6417
rect 23152 6400 23169 6417
rect 23313 6400 23330 6417
rect 24187 6400 24204 6417
rect 24440 6400 24457 6417
rect 24624 6400 24641 6417
rect 28212 6400 28229 6417
rect 28367 6400 28384 6417
rect 6592 6366 6609 6383
rect 7604 6366 7621 6383
rect 29247 6366 29264 6383
rect 16114 6332 16131 6349
rect 6224 6298 6241 6315
rect 6270 6298 6287 6315
rect 16528 6298 16545 6315
rect 6960 6196 6977 6213
rect 5488 6128 5505 6145
rect 5626 6128 5643 6145
rect 6868 6128 6885 6145
rect 7420 6128 7437 6145
rect 20208 6128 20225 6145
rect 6776 6094 6793 6111
rect 6960 6094 6977 6111
rect 7558 6094 7575 6111
rect 7788 6094 7805 6111
rect 11210 6094 11227 6111
rect 19886 6094 19903 6111
rect 20024 6094 20041 6111
rect 20116 6094 20133 6111
rect 6500 6060 6517 6077
rect 7420 6060 7437 6077
rect 7604 6060 7621 6077
rect 6822 6026 6839 6043
rect 7512 6026 7529 6043
rect 11261 6026 11278 6043
rect 11054 5924 11071 5941
rect 29339 5924 29356 5941
rect 9490 5890 9507 5907
rect 10272 5890 10289 5907
rect 10962 5890 10979 5907
rect 18966 5890 18983 5907
rect 20208 5890 20225 5907
rect 26625 5890 26642 5907
rect 28515 5890 28532 5907
rect 7696 5856 7713 5873
rect 7788 5856 7805 5873
rect 8156 5856 8173 5873
rect 9306 5856 9323 5873
rect 9353 5856 9370 5873
rect 9444 5856 9461 5873
rect 9539 5856 9556 5873
rect 9858 5856 9875 5873
rect 9996 5856 10013 5873
rect 10134 5856 10151 5873
rect 10180 5856 10197 5873
rect 11100 5856 11117 5873
rect 11560 5856 11577 5873
rect 17080 5856 17097 5873
rect 17126 5856 17143 5873
rect 17356 5856 17373 5873
rect 18368 5856 18385 5873
rect 18552 5856 18569 5873
rect 18736 5856 18753 5873
rect 19840 5856 19857 5873
rect 20070 5856 20087 5873
rect 26573 5856 26590 5873
rect 28459 5856 28476 5873
rect 8110 5822 8127 5839
rect 11606 5822 11623 5839
rect 11698 5822 11715 5839
rect 20116 5822 20133 5839
rect 26418 5822 26435 5839
rect 28304 5822 28321 5839
rect 9628 5788 9645 5805
rect 10962 5788 10979 5805
rect 7696 5754 7713 5771
rect 8294 5754 8311 5771
rect 11652 5754 11669 5771
rect 17218 5754 17235 5771
rect 27453 5754 27470 5771
rect 10272 5652 10289 5669
rect 17954 5652 17971 5669
rect 18690 5652 18707 5669
rect 19840 5652 19857 5669
rect 7834 5618 7851 5635
rect 7880 5584 7897 5601
rect 10180 5584 10197 5601
rect 10318 5584 10335 5601
rect 16896 5584 16913 5601
rect 16988 5584 17005 5601
rect 26924 5584 26941 5601
rect 7834 5550 7851 5567
rect 7926 5550 7943 5567
rect 8018 5550 8035 5567
rect 8524 5550 8541 5567
rect 8616 5550 8633 5567
rect 8938 5550 8955 5567
rect 9030 5550 9047 5567
rect 9076 5550 9093 5567
rect 10226 5550 10243 5567
rect 15700 5550 15717 5567
rect 15746 5550 15763 5567
rect 16850 5550 16867 5567
rect 17264 5550 17281 5567
rect 18506 5550 18523 5567
rect 18552 5550 18569 5567
rect 18598 5550 18615 5567
rect 19794 5550 19811 5567
rect 20070 5550 20087 5567
rect 22140 5550 22157 5567
rect 22217 5550 22234 5567
rect 22298 5550 22315 5567
rect 22353 5550 22370 5567
rect 22401 5540 22418 5557
rect 22452 5550 22469 5567
rect 26740 5550 26757 5567
rect 26878 5550 26895 5567
rect 27200 5550 27217 5567
rect 27292 5550 27309 5567
rect 7742 5516 7759 5533
rect 8708 5516 8725 5533
rect 15838 5516 15855 5533
rect 17398 5516 17415 5533
rect 27246 5516 27263 5533
rect 9076 5482 9093 5499
rect 15700 5482 15717 5499
rect 16988 5482 17005 5499
rect 22370 5482 22387 5499
rect 7834 5380 7851 5397
rect 9122 5380 9139 5397
rect 10134 5380 10151 5397
rect 15976 5380 15993 5397
rect 16068 5380 16085 5397
rect 17402 5380 17419 5397
rect 22117 5380 22134 5397
rect 25360 5380 25377 5397
rect 15144 5346 15161 5363
rect 20300 5346 20317 5363
rect 21293 5346 21310 5363
rect 24003 5346 24020 5363
rect 7788 5312 7805 5329
rect 7972 5312 7989 5329
rect 8202 5312 8219 5329
rect 8294 5312 8311 5329
rect 8938 5312 8955 5329
rect 8985 5312 9002 5329
rect 10042 5312 10059 5329
rect 10134 5312 10151 5329
rect 15010 5312 15027 5329
rect 15930 5312 15947 5329
rect 16114 5312 16131 5329
rect 17356 5312 17373 5329
rect 17448 5312 17465 5329
rect 18368 5312 18385 5329
rect 19932 5312 19949 5329
rect 20162 5312 20179 5329
rect 21082 5312 21099 5329
rect 21243 5312 21260 5329
rect 23796 5312 23813 5329
rect 23957 5312 23974 5329
rect 25360 5312 25377 5329
rect 25417 5312 25434 5329
rect 25511 5312 25528 5329
rect 25566 5323 25583 5340
rect 25621 5312 25638 5329
rect 25672 5312 25689 5329
rect 7880 5278 7897 5295
rect 16022 5278 16039 5295
rect 18322 5278 18339 5295
rect 18460 5278 18477 5295
rect 24831 5278 24848 5295
rect 7972 5244 7989 5261
rect 8202 5244 8219 5261
rect 15700 5244 15717 5261
rect 18414 5210 18431 5227
rect 8179 5108 8196 5125
rect 22255 5108 22272 5125
rect 25015 5108 25032 5125
rect 18552 5040 18569 5057
rect 19748 5040 19765 5057
rect 21220 5040 21237 5057
rect 23980 5040 23997 5057
rect 8128 5006 8145 5023
rect 18460 5006 18477 5023
rect 18644 5006 18661 5023
rect 19610 5006 19627 5023
rect 19932 5006 19949 5023
rect 21375 5006 21392 5023
rect 24141 5006 24158 5023
rect 21431 4972 21448 4989
rect 24191 4972 24208 4989
rect 18506 4938 18523 4955
rect 18598 4938 18615 4955
rect 16528 4836 16545 4853
rect 19104 4836 19121 4853
rect 16436 4802 16453 4819
rect 17172 4802 17189 4819
rect 18548 4802 18565 4819
rect 21289 4802 21306 4819
rect 22117 4802 22134 4819
rect 16574 4768 16591 4785
rect 17080 4768 17097 4785
rect 17218 4768 17235 4785
rect 19840 4768 19857 4785
rect 20162 4768 20179 4785
rect 21082 4768 21099 4785
rect 21243 4768 21260 4785
rect 18414 4734 18431 4751
rect 19978 4734 19995 4751
rect 16436 4700 16453 4717
rect 17080 4666 17097 4683
rect 17264 4564 17281 4581
rect 25107 4564 25124 4581
rect 16574 4496 16591 4513
rect 24072 4496 24089 4513
rect 16708 4462 16725 4479
rect 24227 4462 24244 4479
rect 24279 4428 24296 4445
rect 18644 3952 18661 3969
rect 19104 3952 19121 3969
rect 18782 3918 18799 3935
<< metal1 >>
rect 3036 29896 29992 29944
rect 15877 29788 15880 29814
rect 15906 29808 15909 29814
rect 15942 29809 15971 29812
rect 15942 29808 15948 29809
rect 15906 29794 15948 29808
rect 15906 29788 15909 29794
rect 15942 29792 15948 29794
rect 15965 29792 15971 29809
rect 15942 29789 15971 29792
rect 15993 29707 16022 29710
rect 15993 29690 15999 29707
rect 16016 29706 16022 29707
rect 16245 29706 16248 29712
rect 16016 29692 16248 29706
rect 16016 29690 16022 29692
rect 15993 29687 16022 29690
rect 16245 29686 16248 29692
rect 16274 29686 16277 29712
rect 3036 29624 29992 29672
rect 10265 29550 10268 29576
rect 10294 29550 10297 29576
rect 11692 29571 11721 29574
rect 11692 29554 11698 29571
rect 11715 29554 11721 29571
rect 11692 29551 11721 29554
rect 11700 29536 11714 29551
rect 15417 29550 15420 29576
rect 15446 29570 15449 29576
rect 15694 29571 15723 29574
rect 15694 29570 15700 29571
rect 15446 29556 15700 29570
rect 15446 29550 15449 29556
rect 15694 29554 15700 29556
rect 15717 29554 15723 29571
rect 15694 29551 15723 29554
rect 16108 29537 16137 29540
rect 16108 29536 16114 29537
rect 11700 29522 12082 29536
rect 10266 29503 10295 29506
rect 10266 29486 10272 29503
rect 10289 29502 10295 29503
rect 10357 29502 10360 29508
rect 10289 29488 10360 29502
rect 10289 29486 10295 29488
rect 10266 29483 10295 29486
rect 10357 29482 10360 29488
rect 10386 29482 10389 29508
rect 10404 29503 10433 29506
rect 10404 29486 10410 29503
rect 10427 29502 10433 29503
rect 10495 29502 10498 29508
rect 10427 29488 10498 29502
rect 10427 29486 10433 29488
rect 10404 29483 10433 29486
rect 10495 29482 10498 29488
rect 10524 29482 10527 29508
rect 11369 29482 11372 29508
rect 11398 29502 11401 29508
rect 12068 29506 12082 29522
rect 15794 29522 16114 29536
rect 11830 29503 11859 29506
rect 11830 29502 11836 29503
rect 11398 29488 11836 29502
rect 11398 29482 11401 29488
rect 11830 29486 11836 29488
rect 11853 29486 11859 29503
rect 11830 29483 11859 29486
rect 12060 29503 12089 29506
rect 12060 29486 12066 29503
rect 12083 29486 12089 29503
rect 12060 29483 12089 29486
rect 12152 29503 12181 29506
rect 12152 29486 12158 29503
rect 12175 29502 12181 29503
rect 12289 29502 12292 29508
rect 12175 29488 12292 29502
rect 12175 29486 12181 29488
rect 12152 29483 12181 29486
rect 12289 29482 12292 29488
rect 12318 29482 12321 29508
rect 15794 29506 15808 29522
rect 16108 29520 16114 29522
rect 16131 29520 16137 29537
rect 16108 29517 16137 29520
rect 16246 29537 16275 29540
rect 16246 29520 16252 29537
rect 16269 29536 16275 29537
rect 16337 29536 16340 29542
rect 16269 29522 16340 29536
rect 16269 29520 16275 29522
rect 16246 29517 16275 29520
rect 16337 29516 16340 29522
rect 16366 29516 16369 29542
rect 15786 29503 15815 29506
rect 15786 29486 15792 29503
rect 15809 29486 15815 29503
rect 15786 29483 15815 29486
rect 15832 29503 15861 29506
rect 15832 29486 15838 29503
rect 15855 29486 15861 29503
rect 15832 29483 15861 29486
rect 16154 29503 16183 29506
rect 16154 29486 16160 29503
rect 16177 29502 16183 29503
rect 16199 29502 16202 29508
rect 16177 29488 16202 29502
rect 16177 29486 16183 29488
rect 16154 29483 16183 29486
rect 8701 29448 8704 29474
rect 8730 29468 8733 29474
rect 11692 29469 11721 29472
rect 8730 29454 11047 29468
rect 8730 29448 8733 29454
rect 10358 29435 10387 29438
rect 10358 29418 10364 29435
rect 10381 29434 10387 29435
rect 10541 29434 10544 29440
rect 10381 29420 10544 29434
rect 10381 29418 10387 29420
rect 10358 29415 10387 29418
rect 10541 29414 10544 29420
rect 10570 29414 10573 29440
rect 11033 29434 11047 29454
rect 11692 29452 11698 29469
rect 11715 29468 11721 29469
rect 11875 29468 11878 29474
rect 11715 29454 11878 29468
rect 11715 29452 11721 29454
rect 11692 29449 11721 29452
rect 11875 29448 11878 29454
rect 11904 29448 11907 29474
rect 12335 29468 12338 29474
rect 11930 29454 12338 29468
rect 11784 29435 11813 29438
rect 11784 29434 11790 29435
rect 11033 29420 11790 29434
rect 11784 29418 11790 29420
rect 11807 29434 11813 29435
rect 11930 29434 11944 29454
rect 12335 29448 12338 29454
rect 12364 29448 12367 29474
rect 15693 29448 15696 29474
rect 15722 29448 15725 29474
rect 15840 29468 15854 29483
rect 16162 29468 16176 29483
rect 16199 29482 16202 29488
rect 16228 29482 16231 29508
rect 15840 29454 16176 29468
rect 11807 29420 11944 29434
rect 11807 29418 11813 29420
rect 11784 29415 11813 29418
rect 12105 29414 12108 29440
rect 12134 29414 12137 29440
rect 15785 29414 15788 29440
rect 15814 29414 15817 29440
rect 16246 29435 16275 29438
rect 16246 29418 16252 29435
rect 16269 29434 16275 29435
rect 16383 29434 16386 29440
rect 16269 29420 16386 29434
rect 16269 29418 16275 29420
rect 16246 29415 16275 29418
rect 16383 29414 16386 29420
rect 16412 29414 16415 29440
rect 3036 29352 29992 29400
rect 14590 29333 14619 29336
rect 14590 29316 14596 29333
rect 14613 29332 14619 29333
rect 15693 29332 15696 29338
rect 14613 29318 15696 29332
rect 14613 29316 14619 29318
rect 14590 29313 14619 29316
rect 15693 29312 15696 29318
rect 15722 29312 15725 29338
rect 15785 29312 15788 29338
rect 15814 29332 15817 29338
rect 16614 29333 16643 29336
rect 16614 29332 16620 29333
rect 15814 29318 16620 29332
rect 15814 29312 15817 29318
rect 16614 29316 16620 29318
rect 16637 29316 16643 29333
rect 16614 29313 16643 29316
rect 7045 29302 7048 29304
rect 7027 29299 7048 29302
rect 7027 29282 7033 29299
rect 7074 29298 7077 29304
rect 10124 29299 10153 29302
rect 7074 29284 7160 29298
rect 7027 29279 7048 29282
rect 7045 29278 7048 29279
rect 7074 29278 7077 29284
rect 6953 29244 6956 29270
rect 6982 29268 6985 29270
rect 6982 29265 7000 29268
rect 6994 29248 7000 29265
rect 7146 29264 7160 29284
rect 10124 29282 10130 29299
rect 10147 29298 10153 29299
rect 10265 29298 10268 29304
rect 10147 29284 10268 29298
rect 10147 29282 10153 29284
rect 10124 29279 10153 29282
rect 10265 29278 10268 29284
rect 10294 29278 10297 29304
rect 11780 29299 11809 29302
rect 11780 29282 11786 29299
rect 11803 29298 11809 29299
rect 12105 29298 12108 29304
rect 11803 29284 12108 29298
rect 11803 29282 11809 29284
rect 11780 29279 11809 29282
rect 12105 29278 12108 29284
rect 12134 29278 12137 29304
rect 15138 29299 15167 29302
rect 14644 29284 15118 29298
rect 8701 29264 8704 29270
rect 7146 29250 8704 29264
rect 6982 29245 7000 29248
rect 6982 29244 6985 29245
rect 8701 29244 8704 29250
rect 8730 29244 8733 29270
rect 8793 29244 8796 29270
rect 8822 29264 8825 29270
rect 8886 29265 8915 29268
rect 8886 29264 8892 29265
rect 8822 29250 8892 29264
rect 8822 29244 8825 29250
rect 8886 29248 8892 29250
rect 8909 29248 8915 29265
rect 8886 29245 8915 29248
rect 8978 29265 9007 29268
rect 8978 29248 8984 29265
rect 9001 29264 9007 29265
rect 9023 29264 9026 29270
rect 9001 29250 9026 29264
rect 9001 29248 9007 29250
rect 8978 29245 9007 29248
rect 9023 29244 9026 29250
rect 9052 29244 9055 29270
rect 9990 29265 10019 29268
rect 9990 29248 9996 29265
rect 10013 29264 10019 29265
rect 10311 29264 10314 29270
rect 10013 29250 10314 29264
rect 10013 29248 10019 29250
rect 9990 29245 10019 29248
rect 10311 29244 10314 29250
rect 10340 29264 10343 29270
rect 11646 29265 11675 29268
rect 11646 29264 11652 29265
rect 10340 29250 11652 29264
rect 10340 29244 10343 29250
rect 11646 29248 11652 29250
rect 11669 29248 11675 29265
rect 11646 29245 11675 29248
rect 13298 29265 13327 29268
rect 13298 29248 13304 29265
rect 13321 29264 13327 29265
rect 13807 29264 13810 29270
rect 13321 29250 13810 29264
rect 13321 29248 13327 29250
rect 13298 29245 13327 29248
rect 13807 29244 13810 29250
rect 13836 29244 13839 29270
rect 14313 29244 14316 29270
rect 14342 29264 14345 29270
rect 14544 29265 14573 29268
rect 14544 29264 14550 29265
rect 14342 29250 14550 29264
rect 14342 29244 14345 29250
rect 14544 29248 14550 29250
rect 14567 29248 14573 29265
rect 14544 29245 14573 29248
rect 6723 29210 6726 29236
rect 6752 29230 6755 29236
rect 6816 29231 6845 29234
rect 6816 29230 6822 29231
rect 6752 29216 6822 29230
rect 6752 29210 6755 29216
rect 6816 29214 6822 29216
rect 6839 29214 6845 29231
rect 6816 29211 6845 29214
rect 13117 29210 13120 29236
rect 13146 29230 13149 29236
rect 14644 29234 14658 29284
rect 14728 29265 14757 29268
rect 14728 29248 14734 29265
rect 14751 29248 14757 29265
rect 15104 29264 15118 29284
rect 15138 29282 15144 29299
rect 15161 29298 15167 29299
rect 15187 29298 15190 29304
rect 15161 29284 15190 29298
rect 15161 29282 15167 29284
rect 15138 29279 15167 29282
rect 15187 29278 15190 29284
rect 15216 29278 15219 29304
rect 15785 29264 15788 29270
rect 15104 29250 15788 29264
rect 14728 29245 14757 29248
rect 13164 29231 13193 29234
rect 13164 29230 13170 29231
rect 13146 29216 13170 29230
rect 13146 29210 13149 29216
rect 13164 29214 13170 29216
rect 13187 29214 13193 29231
rect 13164 29211 13193 29214
rect 14636 29231 14665 29234
rect 14636 29214 14642 29231
rect 14659 29214 14665 29231
rect 14636 29211 14665 29214
rect 13854 29197 13883 29200
rect 13854 29180 13860 29197
rect 13877 29196 13883 29197
rect 13945 29196 13948 29202
rect 13877 29182 13948 29196
rect 13877 29180 13883 29182
rect 13854 29177 13883 29180
rect 13945 29176 13948 29182
rect 13974 29196 13977 29202
rect 14736 29196 14750 29245
rect 15785 29244 15788 29250
rect 15814 29244 15817 29270
rect 16058 29265 16087 29268
rect 16058 29248 16064 29265
rect 16081 29264 16087 29265
rect 16291 29264 16294 29270
rect 16081 29250 16294 29264
rect 16081 29248 16087 29250
rect 16058 29245 16087 29248
rect 16291 29244 16294 29250
rect 16320 29244 16323 29270
rect 15003 29210 15006 29236
rect 15032 29210 15035 29236
rect 15923 29230 15926 29236
rect 15518 29216 15926 29230
rect 13974 29182 14750 29196
rect 13974 29176 13977 29182
rect 7851 29163 7880 29166
rect 7851 29146 7857 29163
rect 7874 29162 7880 29163
rect 8057 29162 8060 29168
rect 7874 29148 8060 29162
rect 7874 29146 7880 29148
rect 7851 29143 7880 29146
rect 8057 29142 8060 29148
rect 8086 29142 8089 29168
rect 8931 29142 8934 29168
rect 8960 29142 8963 29168
rect 10541 29142 10544 29168
rect 10570 29162 10573 29168
rect 10680 29163 10709 29166
rect 10680 29162 10686 29163
rect 10570 29148 10686 29162
rect 10570 29142 10573 29148
rect 10680 29146 10686 29148
rect 10703 29146 10709 29163
rect 10680 29143 10709 29146
rect 11645 29142 11648 29168
rect 11674 29162 11677 29168
rect 12336 29163 12365 29166
rect 12336 29162 12342 29163
rect 11674 29148 12342 29162
rect 11674 29142 11677 29148
rect 12336 29146 12342 29148
rect 12359 29146 12365 29163
rect 12336 29143 12365 29146
rect 13899 29142 13902 29168
rect 13928 29162 13931 29168
rect 14728 29163 14757 29166
rect 14728 29162 14734 29163
rect 13928 29148 14734 29162
rect 13928 29142 13931 29148
rect 14728 29146 14734 29148
rect 14751 29146 14757 29163
rect 14728 29143 14757 29146
rect 15003 29142 15006 29168
rect 15032 29162 15035 29168
rect 15518 29162 15532 29216
rect 15923 29210 15926 29216
rect 15952 29210 15955 29236
rect 15032 29148 15532 29162
rect 15694 29163 15723 29166
rect 15032 29142 15035 29148
rect 15694 29146 15700 29163
rect 15717 29162 15723 29163
rect 15877 29162 15880 29168
rect 15717 29148 15880 29162
rect 15717 29146 15723 29148
rect 15694 29143 15723 29146
rect 15877 29142 15880 29148
rect 15906 29142 15909 29168
rect 3036 29080 29992 29128
rect 6908 29061 6937 29064
rect 6908 29044 6914 29061
rect 6931 29060 6937 29061
rect 6953 29060 6956 29066
rect 6931 29046 6956 29060
rect 6931 29044 6937 29046
rect 6908 29041 6937 29044
rect 6953 29040 6956 29046
rect 6982 29040 6985 29066
rect 10357 29040 10360 29066
rect 10386 29040 10389 29066
rect 11369 29040 11372 29066
rect 11398 29040 11401 29066
rect 11875 29040 11878 29066
rect 11904 29040 11907 29066
rect 13762 29061 13791 29064
rect 13762 29044 13768 29061
rect 13785 29060 13791 29061
rect 13807 29060 13810 29066
rect 13785 29046 13810 29060
rect 13785 29044 13791 29046
rect 13762 29041 13791 29044
rect 13807 29040 13810 29046
rect 13836 29040 13839 29066
rect 15142 29061 15171 29064
rect 15142 29044 15148 29061
rect 15165 29060 15171 29061
rect 15187 29060 15190 29066
rect 15165 29046 15190 29060
rect 15165 29044 15171 29046
rect 15142 29041 15171 29044
rect 15187 29040 15190 29046
rect 15216 29040 15219 29066
rect 16291 29040 16294 29066
rect 16320 29060 16323 29066
rect 16384 29061 16413 29064
rect 16384 29060 16390 29061
rect 16320 29046 16390 29060
rect 16320 29040 16323 29046
rect 16384 29044 16390 29046
rect 16407 29044 16413 29061
rect 16384 29041 16413 29044
rect 8655 29006 8658 29032
rect 8684 29026 8687 29032
rect 8817 29027 8846 29030
rect 8817 29026 8823 29027
rect 8684 29012 8823 29026
rect 8684 29006 8687 29012
rect 8817 29010 8823 29012
rect 8840 29010 8846 29027
rect 8817 29007 8846 29010
rect 8885 29006 8888 29032
rect 8914 29026 8917 29032
rect 8914 29012 9046 29026
rect 8914 29006 8917 29012
rect 8388 28978 9000 28992
rect 4699 28938 4702 28964
rect 4728 28958 4731 28964
rect 6815 28962 6818 28964
rect 4792 28959 4821 28962
rect 4792 28958 4798 28959
rect 4728 28944 4798 28958
rect 4728 28938 4731 28944
rect 4792 28942 4798 28944
rect 4815 28942 4821 28959
rect 4792 28939 4821 28942
rect 6724 28959 6753 28962
rect 6724 28942 6730 28959
rect 6747 28942 6753 28959
rect 6724 28939 6753 28942
rect 6793 28959 6818 28962
rect 6793 28942 6799 28959
rect 6816 28942 6818 28959
rect 6793 28939 6818 28942
rect 4929 28904 4932 28930
rect 4958 28904 4961 28930
rect 5573 28924 5576 28930
rect 5543 28910 5576 28924
rect 5573 28904 5576 28910
rect 5602 28904 5605 28930
rect 6732 28924 6746 28939
rect 6815 28938 6818 28939
rect 6844 28938 6847 28964
rect 6861 28938 6864 28964
rect 6890 28938 6893 28964
rect 6954 28959 6983 28962
rect 6954 28942 6960 28959
rect 6977 28958 6983 28959
rect 7414 28959 7443 28962
rect 6977 28944 7390 28958
rect 6977 28942 6983 28944
rect 6954 28939 6983 28942
rect 7321 28924 7324 28930
rect 6732 28910 7324 28924
rect 7321 28904 7324 28910
rect 7350 28904 7353 28930
rect 5619 28870 5622 28896
rect 5648 28890 5651 28896
rect 5666 28891 5695 28894
rect 5666 28890 5672 28891
rect 5648 28876 5672 28890
rect 5648 28870 5651 28876
rect 5666 28874 5672 28876
rect 5689 28874 5695 28891
rect 7376 28890 7390 28944
rect 7414 28942 7420 28959
rect 7437 28942 7443 28959
rect 7414 28939 7443 28942
rect 7422 28924 7436 28939
rect 7459 28938 7462 28964
rect 7488 28938 7491 28964
rect 7505 28938 7508 28964
rect 7534 28938 7537 28964
rect 8057 28938 8060 28964
rect 8086 28958 8089 28964
rect 8388 28958 8402 28978
rect 8086 28944 8402 28958
rect 8086 28938 8089 28944
rect 8425 28938 8428 28964
rect 8454 28938 8457 28964
rect 8518 28959 8547 28962
rect 8518 28942 8524 28959
rect 8541 28958 8547 28959
rect 8748 28959 8777 28962
rect 8748 28958 8754 28959
rect 8541 28944 8754 28958
rect 8541 28942 8547 28944
rect 8518 28939 8547 28942
rect 8748 28942 8754 28944
rect 8771 28942 8777 28959
rect 8748 28939 8777 28942
rect 8886 28959 8915 28962
rect 8886 28942 8892 28959
rect 8909 28958 8915 28959
rect 8931 28958 8934 28964
rect 8909 28944 8934 28958
rect 8909 28942 8915 28944
rect 8886 28939 8915 28942
rect 8149 28924 8152 28930
rect 7422 28910 8152 28924
rect 8149 28904 8152 28910
rect 8178 28924 8181 28930
rect 8472 28925 8501 28928
rect 8472 28924 8478 28925
rect 8178 28910 8478 28924
rect 8178 28904 8181 28910
rect 8472 28908 8478 28910
rect 8495 28908 8501 28925
rect 8756 28924 8770 28939
rect 8931 28938 8934 28944
rect 8960 28938 8963 28964
rect 8986 28962 9000 28978
rect 8978 28959 9007 28962
rect 8978 28942 8984 28959
rect 9001 28942 9007 28959
rect 9032 28958 9046 29012
rect 13117 29006 13120 29032
rect 13146 29026 13149 29032
rect 15003 29026 15006 29032
rect 13146 29012 15006 29026
rect 13146 29006 13149 29012
rect 15003 29006 15006 29012
rect 15032 29006 15035 29032
rect 15693 29006 15696 29032
rect 15722 29006 15725 29032
rect 10403 28972 10406 28998
rect 10432 28972 10435 28998
rect 10541 28972 10544 28998
rect 10570 28992 10573 28998
rect 11140 28993 11169 28996
rect 11140 28992 11146 28993
rect 10570 28978 11146 28992
rect 10570 28972 10573 28978
rect 11140 28976 11146 28978
rect 11163 28976 11169 28993
rect 13899 28992 13902 28998
rect 11140 28973 11169 28976
rect 13816 28978 13902 28992
rect 10266 28959 10295 28962
rect 10266 28958 10272 28959
rect 9032 28944 10272 28958
rect 8978 28939 9007 28942
rect 10266 28942 10272 28944
rect 10289 28942 10295 28959
rect 10266 28939 10295 28942
rect 10312 28959 10341 28962
rect 10312 28942 10318 28959
rect 10335 28958 10341 28959
rect 10495 28958 10498 28964
rect 10335 28944 10498 28958
rect 10335 28942 10341 28944
rect 10312 28939 10341 28942
rect 9299 28924 9302 28930
rect 8756 28910 9302 28924
rect 8472 28905 8501 28908
rect 9299 28904 9302 28910
rect 9328 28904 9331 28930
rect 10274 28924 10288 28939
rect 10495 28938 10498 28944
rect 10524 28938 10527 28964
rect 11185 28938 11188 28964
rect 11214 28958 11217 28964
rect 11645 28958 11648 28964
rect 11214 28944 11648 28958
rect 11214 28938 11217 28944
rect 11645 28938 11648 28944
rect 11674 28958 11677 28964
rect 11692 28959 11721 28962
rect 11692 28958 11698 28959
rect 11674 28944 11698 28958
rect 11674 28938 11677 28944
rect 11692 28942 11698 28944
rect 11715 28942 11721 28959
rect 11692 28939 11721 28942
rect 11783 28938 11786 28964
rect 11812 28938 11815 28964
rect 13762 28959 13791 28962
rect 13762 28942 13768 28959
rect 13785 28958 13791 28959
rect 13816 28958 13830 28978
rect 13899 28972 13902 28978
rect 13928 28972 13931 28998
rect 15417 28992 15420 28998
rect 15196 28978 15420 28992
rect 13785 28944 13830 28958
rect 13854 28959 13883 28962
rect 13785 28942 13791 28944
rect 13762 28939 13791 28942
rect 13854 28942 13860 28959
rect 13877 28942 13883 28959
rect 13854 28939 13883 28942
rect 10357 28924 10360 28930
rect 10274 28910 10360 28924
rect 10357 28904 10360 28910
rect 10386 28924 10389 28930
rect 10541 28924 10544 28930
rect 10386 28910 10544 28924
rect 10386 28904 10389 28910
rect 10541 28904 10544 28910
rect 10570 28904 10573 28930
rect 13862 28924 13876 28939
rect 14083 28938 14086 28964
rect 14112 28962 14115 28964
rect 14112 28959 14131 28962
rect 14125 28942 14131 28959
rect 14112 28939 14131 28942
rect 15142 28959 15171 28962
rect 15142 28942 15148 28959
rect 15165 28958 15171 28959
rect 15196 28958 15210 28978
rect 15417 28972 15420 28978
rect 15446 28972 15449 28998
rect 16292 28993 16321 28996
rect 16292 28992 16298 28993
rect 15794 28978 16298 28992
rect 15794 28964 15808 28978
rect 16292 28976 16298 28978
rect 16315 28976 16321 28993
rect 16292 28973 16321 28976
rect 17082 28978 17188 28992
rect 17082 28964 17096 28978
rect 15165 28944 15210 28958
rect 15234 28959 15263 28962
rect 15165 28942 15171 28944
rect 15142 28939 15171 28942
rect 15234 28942 15240 28959
rect 15257 28942 15263 28959
rect 15234 28939 15263 28942
rect 14112 28938 14115 28939
rect 13862 28910 14382 28924
rect 8932 28891 8961 28894
rect 8932 28890 8938 28891
rect 7376 28876 8938 28890
rect 5666 28871 5695 28874
rect 8932 28874 8938 28876
rect 8955 28874 8961 28891
rect 8932 28871 8961 28874
rect 14153 28891 14182 28894
rect 14153 28874 14159 28891
rect 14176 28890 14182 28891
rect 14313 28890 14316 28896
rect 14176 28876 14316 28890
rect 14176 28874 14182 28876
rect 14153 28871 14182 28874
rect 14313 28870 14316 28876
rect 14342 28870 14345 28896
rect 14368 28890 14382 28910
rect 14589 28890 14592 28896
rect 14368 28876 14592 28890
rect 14589 28870 14592 28876
rect 14618 28890 14621 28896
rect 15242 28890 15256 28939
rect 15785 28938 15788 28964
rect 15814 28938 15817 28964
rect 15832 28959 15861 28962
rect 15832 28942 15838 28959
rect 15855 28958 15861 28959
rect 15877 28958 15880 28964
rect 15855 28944 15880 28958
rect 15855 28942 15861 28944
rect 15832 28939 15861 28942
rect 15877 28938 15880 28944
rect 15906 28938 15909 28964
rect 16199 28938 16202 28964
rect 16228 28938 16231 28964
rect 16245 28938 16248 28964
rect 16274 28938 16277 28964
rect 16383 28938 16386 28964
rect 16412 28938 16415 28964
rect 17027 28938 17030 28964
rect 17056 28938 17059 28964
rect 17073 28938 17076 28964
rect 17102 28938 17105 28964
rect 17120 28959 17149 28962
rect 17120 28942 17126 28959
rect 17143 28942 17149 28959
rect 17174 28958 17188 28978
rect 17442 28959 17471 28962
rect 17442 28958 17448 28959
rect 17174 28944 17448 28958
rect 17120 28939 17149 28942
rect 17442 28942 17448 28944
rect 17465 28942 17471 28959
rect 17442 28939 17471 28942
rect 17534 28959 17563 28962
rect 17534 28942 17540 28959
rect 17557 28942 17563 28959
rect 17534 28939 17563 28942
rect 15694 28925 15723 28928
rect 15694 28908 15700 28925
rect 15717 28924 15723 28925
rect 15739 28924 15742 28930
rect 15717 28910 15742 28924
rect 15717 28908 15723 28910
rect 15694 28905 15723 28908
rect 15739 28904 15742 28910
rect 15768 28904 15771 28930
rect 17128 28924 17142 28939
rect 17165 28924 17168 28930
rect 17128 28910 17168 28924
rect 17165 28904 17168 28910
rect 17194 28924 17197 28930
rect 17542 28924 17556 28939
rect 17194 28910 17556 28924
rect 17626 28925 17655 28928
rect 17194 28904 17197 28910
rect 17626 28908 17632 28925
rect 17649 28924 17655 28925
rect 17671 28924 17674 28930
rect 17649 28910 17674 28924
rect 17649 28908 17655 28910
rect 17626 28905 17655 28908
rect 17671 28904 17674 28910
rect 17700 28904 17703 28930
rect 14618 28876 15256 28890
rect 14618 28870 14621 28876
rect 17211 28870 17214 28896
rect 17240 28870 17243 28896
rect 3036 28808 29992 28856
rect 5527 28768 5530 28794
rect 5556 28788 5559 28794
rect 5574 28789 5603 28792
rect 5574 28788 5580 28789
rect 5556 28774 5580 28788
rect 5556 28768 5559 28774
rect 5574 28772 5580 28774
rect 5597 28772 5603 28789
rect 5574 28769 5603 28772
rect 6815 28768 6818 28794
rect 6844 28788 6847 28794
rect 6908 28789 6937 28792
rect 6908 28788 6914 28789
rect 6844 28774 6914 28788
rect 6844 28768 6847 28774
rect 6908 28772 6914 28774
rect 6931 28772 6937 28789
rect 6908 28769 6937 28772
rect 6953 28768 6956 28794
rect 6982 28788 6985 28794
rect 8379 28788 8382 28794
rect 6982 28774 8382 28788
rect 6982 28768 6985 28774
rect 8379 28768 8382 28774
rect 8408 28768 8411 28794
rect 8425 28768 8428 28794
rect 8454 28788 8457 28794
rect 8840 28789 8869 28792
rect 8840 28788 8846 28789
rect 8454 28774 8846 28788
rect 8454 28768 8457 28774
rect 8840 28772 8846 28774
rect 8863 28772 8869 28789
rect 8840 28769 8869 28772
rect 15832 28789 15861 28792
rect 15832 28772 15838 28789
rect 15855 28788 15861 28789
rect 16199 28788 16202 28794
rect 15855 28774 16202 28788
rect 15855 28772 15861 28774
rect 15832 28769 15861 28772
rect 16199 28768 16202 28774
rect 16228 28768 16231 28794
rect 17027 28768 17030 28794
rect 17056 28788 17059 28794
rect 18085 28788 18088 28794
rect 17056 28774 18088 28788
rect 17056 28768 17059 28774
rect 18085 28768 18088 28774
rect 18114 28788 18117 28794
rect 18114 28774 18476 28788
rect 18114 28768 18117 28774
rect 5987 28754 5990 28760
rect 5451 28740 5990 28754
rect 5582 28726 5596 28740
rect 5987 28734 5990 28740
rect 6016 28754 6019 28760
rect 6264 28755 6293 28758
rect 6264 28754 6270 28755
rect 6016 28740 6270 28754
rect 6016 28734 6019 28740
rect 6264 28738 6270 28740
rect 6287 28738 6293 28755
rect 6264 28735 6293 28738
rect 6677 28734 6680 28760
rect 6706 28754 6709 28760
rect 7505 28754 7508 28760
rect 6706 28740 7508 28754
rect 6706 28734 6709 28740
rect 7505 28734 7508 28740
rect 7534 28754 7537 28760
rect 8655 28754 8658 28760
rect 7534 28740 8658 28754
rect 7534 28734 7537 28740
rect 5573 28700 5576 28726
rect 5602 28700 5605 28726
rect 6585 28700 6588 28726
rect 6614 28700 6617 28726
rect 6815 28700 6818 28726
rect 6844 28720 6847 28726
rect 6862 28721 6891 28724
rect 6862 28720 6868 28721
rect 6844 28706 6868 28720
rect 6844 28700 6847 28706
rect 6862 28704 6868 28706
rect 6885 28704 6891 28721
rect 6862 28701 6891 28704
rect 6953 28700 6956 28726
rect 6982 28700 6985 28726
rect 7000 28721 7029 28724
rect 7000 28704 7006 28721
rect 7023 28720 7029 28721
rect 7689 28720 7692 28726
rect 7023 28706 7692 28720
rect 7023 28704 7029 28706
rect 7000 28701 7029 28704
rect 7689 28700 7692 28706
rect 7718 28700 7721 28726
rect 8112 28724 8126 28740
rect 8655 28734 8658 28740
rect 8684 28734 8687 28760
rect 10312 28755 10341 28758
rect 10312 28738 10318 28755
rect 10335 28754 10341 28755
rect 10495 28754 10498 28760
rect 10335 28740 10498 28754
rect 10335 28738 10341 28740
rect 10312 28735 10341 28738
rect 10495 28734 10498 28740
rect 10524 28734 10527 28760
rect 14911 28734 14914 28760
rect 14940 28754 14943 28760
rect 18462 28758 18476 28774
rect 20937 28768 20940 28794
rect 20966 28788 20969 28794
rect 21030 28789 21059 28792
rect 21030 28788 21036 28789
rect 20966 28774 21036 28788
rect 20966 28768 20969 28774
rect 21030 28772 21036 28774
rect 21053 28772 21059 28789
rect 21030 28769 21059 28772
rect 18454 28755 18483 28758
rect 14940 28740 17825 28754
rect 14940 28734 14943 28740
rect 18454 28738 18460 28755
rect 18477 28738 18483 28755
rect 18454 28735 18483 28738
rect 19980 28740 20539 28754
rect 8104 28721 8133 28724
rect 8104 28704 8110 28721
rect 8127 28704 8133 28721
rect 8104 28701 8133 28704
rect 8149 28700 8152 28726
rect 8178 28724 8181 28726
rect 8178 28721 8202 28724
rect 8178 28704 8179 28721
rect 8196 28704 8202 28721
rect 8178 28701 8202 28704
rect 8334 28721 8363 28724
rect 8334 28704 8340 28721
rect 8357 28704 8363 28721
rect 8334 28701 8363 28704
rect 8178 28700 8181 28701
rect 4699 28666 4702 28692
rect 4728 28666 4731 28692
rect 4838 28687 4867 28690
rect 4838 28670 4844 28687
rect 4861 28686 4867 28687
rect 5159 28686 5162 28692
rect 4861 28672 5162 28686
rect 4861 28670 4867 28672
rect 4838 28667 4867 28670
rect 5159 28666 5162 28672
rect 5188 28666 5191 28692
rect 6632 28687 6661 28690
rect 6632 28670 6638 28687
rect 6655 28686 6661 28687
rect 8342 28686 8356 28701
rect 8379 28700 8382 28726
rect 8408 28720 8411 28726
rect 8793 28720 8796 28726
rect 8408 28706 8796 28720
rect 8408 28700 8411 28706
rect 8793 28700 8796 28706
rect 8822 28700 8825 28726
rect 8886 28721 8915 28724
rect 8886 28704 8892 28721
rect 8909 28720 8915 28721
rect 9023 28720 9026 28726
rect 8909 28706 9026 28720
rect 8909 28704 8915 28706
rect 8886 28701 8915 28704
rect 9023 28700 9026 28706
rect 9052 28700 9055 28726
rect 10357 28700 10360 28726
rect 10386 28720 10389 28726
rect 10404 28721 10433 28724
rect 10404 28720 10410 28721
rect 10386 28706 10410 28720
rect 10386 28700 10389 28706
rect 10404 28704 10410 28706
rect 10427 28704 10433 28721
rect 10404 28701 10433 28704
rect 10450 28721 10479 28724
rect 10450 28704 10456 28721
rect 10473 28720 10479 28721
rect 11185 28720 11188 28726
rect 10473 28706 11188 28720
rect 10473 28704 10479 28706
rect 10450 28701 10479 28704
rect 8977 28686 8980 28692
rect 6655 28672 8310 28686
rect 8342 28672 8980 28686
rect 6655 28670 6661 28672
rect 6632 28667 6661 28670
rect 7000 28653 7029 28656
rect 7000 28636 7006 28653
rect 7023 28652 7029 28653
rect 8242 28653 8271 28656
rect 8242 28652 8248 28653
rect 7023 28638 8248 28652
rect 7023 28636 7029 28638
rect 7000 28633 7029 28636
rect 8242 28636 8248 28638
rect 8265 28636 8271 28653
rect 8296 28652 8310 28672
rect 8977 28666 8980 28672
rect 9006 28666 9009 28692
rect 9032 28686 9046 28700
rect 9345 28686 9348 28692
rect 9032 28672 9348 28686
rect 9345 28666 9348 28672
rect 9374 28686 9377 28692
rect 10458 28686 10472 28701
rect 11185 28700 11188 28706
rect 11214 28700 11217 28726
rect 13348 28721 13377 28724
rect 13348 28704 13354 28721
rect 13371 28720 13377 28721
rect 14359 28720 14362 28726
rect 13371 28706 14362 28720
rect 13371 28704 13377 28706
rect 13348 28701 13377 28704
rect 14359 28700 14362 28706
rect 14388 28700 14391 28726
rect 15739 28700 15742 28726
rect 15768 28720 15771 28726
rect 15786 28721 15815 28724
rect 15786 28720 15792 28721
rect 15768 28706 15792 28720
rect 15768 28700 15771 28706
rect 15786 28704 15792 28706
rect 15809 28704 15815 28721
rect 15786 28701 15815 28704
rect 9374 28672 10472 28686
rect 9374 28666 9377 28672
rect 13255 28666 13258 28692
rect 13284 28686 13287 28692
rect 13394 28687 13423 28690
rect 13394 28686 13400 28687
rect 13284 28672 13400 28686
rect 13284 28666 13287 28672
rect 13394 28670 13400 28672
rect 13417 28670 13423 28687
rect 13394 28667 13423 28670
rect 13486 28687 13515 28690
rect 13486 28670 13492 28687
rect 13509 28686 13515 28687
rect 14083 28686 14086 28692
rect 13509 28672 14086 28686
rect 13509 28670 13515 28672
rect 13486 28667 13515 28670
rect 13209 28652 13212 28658
rect 8296 28638 13212 28652
rect 8242 28633 8271 28636
rect 13209 28632 13212 28638
rect 13238 28632 13241 28658
rect 13402 28652 13416 28667
rect 14083 28666 14086 28672
rect 14112 28686 14115 28692
rect 15794 28686 15808 28701
rect 15877 28700 15880 28726
rect 15906 28700 15909 28726
rect 17120 28721 17149 28724
rect 17120 28704 17126 28721
rect 17143 28720 17149 28721
rect 17395 28720 17398 28726
rect 17143 28706 17398 28720
rect 17143 28704 17149 28706
rect 17120 28701 17149 28704
rect 17395 28700 17398 28706
rect 17424 28700 17427 28726
rect 19980 28720 19994 28740
rect 18147 28706 19994 28720
rect 20845 28700 20848 28726
rect 20874 28700 20877 28726
rect 14112 28672 15808 28686
rect 17074 28687 17103 28690
rect 14112 28666 14115 28672
rect 17074 28670 17080 28687
rect 17097 28670 17103 28687
rect 17074 28667 17103 28670
rect 16337 28652 16340 28658
rect 13402 28638 16340 28652
rect 16337 28632 16340 28638
rect 16366 28652 16369 28658
rect 16843 28652 16846 28658
rect 16366 28638 16846 28652
rect 16366 28632 16369 28638
rect 16843 28632 16846 28638
rect 16872 28632 16875 28658
rect 17082 28652 17096 28667
rect 17211 28666 17214 28692
rect 17240 28666 17243 28692
rect 17441 28666 17444 28692
rect 17470 28666 17473 28692
rect 17579 28666 17582 28692
rect 17608 28666 17611 28692
rect 20155 28666 20158 28692
rect 20184 28666 20187 28692
rect 20293 28666 20296 28692
rect 20322 28666 20325 28692
rect 17082 28638 17326 28652
rect 8287 28598 8290 28624
rect 8316 28598 8319 28624
rect 10357 28598 10360 28624
rect 10386 28598 10389 28624
rect 13301 28598 13304 28624
rect 13330 28618 13333 28624
rect 13440 28619 13469 28622
rect 13440 28618 13446 28619
rect 13330 28604 13446 28618
rect 13330 28598 13333 28604
rect 13440 28602 13446 28604
rect 13463 28602 13469 28619
rect 13440 28599 13469 28602
rect 17166 28619 17195 28622
rect 17166 28602 17172 28619
rect 17189 28618 17195 28619
rect 17257 28618 17260 28624
rect 17189 28604 17260 28618
rect 17189 28602 17195 28604
rect 17166 28599 17195 28602
rect 17257 28598 17260 28604
rect 17286 28598 17289 28624
rect 17312 28618 17326 28638
rect 17671 28618 17674 28624
rect 17312 28604 17674 28618
rect 17671 28598 17674 28604
rect 17700 28598 17703 28624
rect 3036 28536 29992 28584
rect 5159 28496 5162 28522
rect 5188 28496 5191 28522
rect 6203 28502 17947 28516
rect 5481 28428 5484 28454
rect 5510 28448 5513 28454
rect 6203 28448 6217 28502
rect 6861 28462 6864 28488
rect 6890 28462 6893 28488
rect 16660 28483 16689 28486
rect 16660 28482 16666 28483
rect 14184 28468 14290 28482
rect 5510 28434 6217 28448
rect 12934 28449 12963 28452
rect 5510 28428 5513 28434
rect 12934 28432 12940 28449
rect 12957 28448 12963 28449
rect 13946 28449 13975 28452
rect 12957 28434 13692 28448
rect 12957 28432 12963 28434
rect 12934 28429 12963 28432
rect 5344 28415 5373 28418
rect 5344 28398 5350 28415
rect 5367 28414 5373 28415
rect 5527 28414 5530 28420
rect 5367 28400 5530 28414
rect 5367 28398 5373 28400
rect 5344 28395 5373 28398
rect 5527 28394 5530 28400
rect 5556 28394 5559 28420
rect 6677 28394 6680 28420
rect 6706 28394 6709 28420
rect 6769 28394 6772 28420
rect 6798 28394 6801 28420
rect 8426 28415 8455 28418
rect 8426 28398 8432 28415
rect 8449 28414 8455 28415
rect 10174 28415 10203 28418
rect 10174 28414 10180 28415
rect 8449 28400 10180 28414
rect 8449 28398 8455 28400
rect 8426 28395 8455 28398
rect 10174 28398 10180 28400
rect 10197 28414 10203 28415
rect 10219 28414 10222 28420
rect 10197 28400 10222 28414
rect 10197 28398 10203 28400
rect 10174 28395 10203 28398
rect 10219 28394 10222 28400
rect 10248 28394 10251 28420
rect 8287 28360 8290 28386
rect 8316 28380 8319 28386
rect 8586 28381 8615 28384
rect 8586 28380 8592 28381
rect 8316 28366 8592 28380
rect 8316 28360 8319 28366
rect 8586 28364 8592 28366
rect 8609 28364 8615 28381
rect 8586 28361 8615 28364
rect 8637 28381 8666 28384
rect 8637 28364 8643 28381
rect 8660 28380 8666 28381
rect 8701 28380 8704 28386
rect 8660 28366 8704 28380
rect 8660 28364 8666 28366
rect 8637 28361 8666 28364
rect 8701 28360 8704 28366
rect 8730 28360 8733 28386
rect 10127 28360 10130 28386
rect 10156 28380 10159 28386
rect 10297 28381 10326 28384
rect 10297 28380 10303 28381
rect 10156 28366 10303 28380
rect 10156 28360 10159 28366
rect 10297 28364 10303 28366
rect 10320 28364 10326 28381
rect 10297 28361 10326 28364
rect 5390 28347 5419 28350
rect 5390 28330 5396 28347
rect 5413 28346 5419 28347
rect 5527 28346 5530 28352
rect 5413 28332 5530 28346
rect 5413 28330 5419 28332
rect 5390 28327 5419 28330
rect 5527 28326 5530 28332
rect 5556 28326 5559 28352
rect 9115 28326 9118 28352
rect 9144 28346 9147 28352
rect 9461 28347 9490 28350
rect 9461 28346 9467 28347
rect 9144 28332 9467 28346
rect 9144 28326 9147 28332
rect 9461 28330 9467 28332
rect 9484 28330 9490 28347
rect 9461 28327 9490 28330
rect 10863 28326 10866 28352
rect 10892 28326 10895 28352
rect 12942 28346 12956 28429
rect 13678 28414 13692 28434
rect 13946 28432 13952 28449
rect 13969 28448 13975 28449
rect 14184 28448 14198 28468
rect 13969 28434 14198 28448
rect 14276 28448 14290 28468
rect 15702 28468 16666 28482
rect 15234 28449 15263 28452
rect 14276 28434 15210 28448
rect 13969 28432 13975 28434
rect 13946 28429 13975 28432
rect 14222 28415 14251 28418
rect 14222 28414 14228 28415
rect 13678 28400 14228 28414
rect 14222 28398 14228 28400
rect 14245 28398 14251 28415
rect 14222 28395 14251 28398
rect 14911 28394 14914 28420
rect 14940 28394 14943 28420
rect 15196 28414 15210 28434
rect 15234 28432 15240 28449
rect 15257 28448 15263 28449
rect 15463 28448 15466 28454
rect 15257 28434 15466 28448
rect 15257 28432 15263 28434
rect 15234 28429 15263 28432
rect 15463 28428 15466 28434
rect 15492 28448 15495 28454
rect 15702 28452 15716 28468
rect 16660 28466 16666 28468
rect 16683 28482 16689 28483
rect 17165 28482 17168 28488
rect 16683 28468 17168 28482
rect 16683 28466 16689 28468
rect 16660 28463 16689 28466
rect 17165 28462 17168 28468
rect 17194 28462 17197 28488
rect 15694 28449 15723 28452
rect 15694 28448 15700 28449
rect 15492 28434 15700 28448
rect 15492 28428 15495 28434
rect 15694 28432 15700 28434
rect 15717 28432 15723 28449
rect 15694 28429 15723 28432
rect 15739 28428 15742 28454
rect 15768 28448 15771 28454
rect 15786 28449 15815 28452
rect 15786 28448 15792 28449
rect 15768 28434 15792 28448
rect 15768 28428 15771 28434
rect 15786 28432 15792 28434
rect 15809 28432 15815 28449
rect 15786 28429 15815 28432
rect 15924 28449 15953 28452
rect 15924 28432 15930 28449
rect 15947 28432 15953 28449
rect 15924 28429 15953 28432
rect 15831 28414 15834 28420
rect 15196 28400 15834 28414
rect 15831 28394 15834 28400
rect 15860 28414 15863 28420
rect 15932 28414 15946 28429
rect 15969 28428 15972 28454
rect 15998 28448 16001 28454
rect 17027 28448 17030 28454
rect 15998 28434 17030 28448
rect 15998 28428 16001 28434
rect 16622 28418 16636 28434
rect 17027 28428 17030 28434
rect 17056 28428 17059 28454
rect 15860 28400 15946 28414
rect 15860 28394 15863 28400
rect 13071 28360 13074 28386
rect 13100 28360 13103 28386
rect 13209 28360 13212 28386
rect 13238 28380 13241 28386
rect 14360 28381 14389 28384
rect 13238 28366 13317 28380
rect 13685 28366 13922 28380
rect 13238 28360 13241 28366
rect 13117 28346 13120 28352
rect 12942 28332 13120 28346
rect 13117 28326 13120 28332
rect 13146 28326 13149 28352
rect 13908 28346 13922 28366
rect 14360 28364 14366 28381
rect 14383 28380 14389 28381
rect 14497 28380 14500 28386
rect 14383 28366 14500 28380
rect 14383 28364 14389 28366
rect 14360 28361 14389 28364
rect 14497 28360 14500 28366
rect 14526 28360 14529 28386
rect 15932 28380 15946 28400
rect 16614 28415 16643 28418
rect 16614 28398 16620 28415
rect 16637 28398 16643 28415
rect 16705 28414 16708 28420
rect 16734 28418 16737 28420
rect 16734 28415 16751 28418
rect 16614 28395 16643 28398
rect 16668 28400 16708 28414
rect 16668 28380 16682 28400
rect 16705 28394 16708 28400
rect 16745 28398 16751 28415
rect 16734 28395 16751 28398
rect 17212 28415 17241 28418
rect 17212 28398 17218 28415
rect 17235 28398 17241 28415
rect 17212 28395 17241 28398
rect 16734 28394 16737 28395
rect 17220 28380 17234 28395
rect 17257 28394 17260 28420
rect 17286 28414 17289 28420
rect 17340 28415 17369 28418
rect 17340 28414 17346 28415
rect 17286 28400 17346 28414
rect 17286 28394 17289 28400
rect 17340 28398 17346 28400
rect 17363 28398 17369 28415
rect 17933 28414 17947 28502
rect 20293 28496 20296 28522
rect 20322 28496 20325 28522
rect 19235 28428 19238 28454
rect 19264 28448 19267 28454
rect 20570 28449 20599 28452
rect 20570 28448 20576 28449
rect 19264 28434 19718 28448
rect 19264 28428 19267 28434
rect 19282 28415 19311 28418
rect 17933 28400 19258 28414
rect 17340 28395 17369 28398
rect 17441 28380 17444 28386
rect 14552 28366 14605 28380
rect 15932 28366 16682 28380
rect 16806 28366 17444 28380
rect 14552 28346 14566 28366
rect 13908 28332 14566 28346
rect 15923 28326 15926 28352
rect 15952 28346 15955 28352
rect 16806 28346 16820 28366
rect 17441 28360 17444 28366
rect 17470 28360 17473 28386
rect 18499 28380 18502 28386
rect 17496 28366 18502 28380
rect 15952 28332 16820 28346
rect 15952 28326 15955 28332
rect 16843 28326 16846 28352
rect 16872 28346 16875 28352
rect 17496 28346 17510 28366
rect 18499 28360 18502 28366
rect 18528 28360 18531 28386
rect 16872 28332 17510 28346
rect 16872 28326 16875 28332
rect 17901 28326 17904 28352
rect 17930 28326 17933 28352
rect 19244 28346 19258 28400
rect 19282 28398 19288 28415
rect 19305 28414 19311 28415
rect 19373 28414 19376 28420
rect 19305 28400 19376 28414
rect 19305 28398 19311 28400
rect 19282 28395 19311 28398
rect 19373 28394 19376 28400
rect 19402 28394 19405 28420
rect 19704 28418 19718 28434
rect 19796 28434 20576 28448
rect 19696 28415 19725 28418
rect 19696 28398 19702 28415
rect 19719 28398 19725 28415
rect 19696 28395 19725 28398
rect 19466 28381 19495 28384
rect 19466 28364 19472 28381
rect 19489 28380 19495 28381
rect 19796 28380 19810 28434
rect 20570 28432 20576 28434
rect 20593 28448 20599 28449
rect 20615 28448 20618 28454
rect 20593 28434 20618 28448
rect 20593 28432 20599 28434
rect 20570 28429 20599 28432
rect 20615 28428 20618 28434
rect 20644 28428 20647 28454
rect 20478 28415 20507 28418
rect 20478 28398 20484 28415
rect 20501 28414 20507 28415
rect 20891 28414 20894 28420
rect 20501 28400 20894 28414
rect 20501 28398 20507 28400
rect 20478 28395 20507 28398
rect 20891 28394 20894 28400
rect 20920 28394 20923 28420
rect 19489 28366 19810 28380
rect 19489 28364 19495 28366
rect 19466 28361 19495 28364
rect 19282 28347 19311 28350
rect 19282 28346 19288 28347
rect 19244 28332 19288 28346
rect 19282 28330 19288 28332
rect 19305 28330 19311 28347
rect 19282 28327 19311 28330
rect 20523 28326 20526 28352
rect 20552 28326 20555 28352
rect 3036 28264 29992 28312
rect 4929 28224 4932 28250
rect 4958 28244 4961 28250
rect 5206 28245 5235 28248
rect 5206 28244 5212 28245
rect 4958 28230 5212 28244
rect 4958 28224 4961 28230
rect 5206 28228 5212 28230
rect 5229 28228 5235 28245
rect 5206 28225 5235 28228
rect 5390 28245 5419 28248
rect 5390 28228 5396 28245
rect 5413 28244 5419 28245
rect 5619 28244 5622 28250
rect 5413 28230 5622 28244
rect 5413 28228 5419 28230
rect 5390 28225 5419 28228
rect 5619 28224 5622 28230
rect 5648 28224 5651 28250
rect 8977 28224 8980 28250
rect 9006 28224 9009 28250
rect 10541 28224 10544 28250
rect 10570 28224 10573 28250
rect 10588 28245 10617 28248
rect 10588 28228 10594 28245
rect 10611 28244 10617 28245
rect 11185 28244 11188 28250
rect 10611 28230 11188 28244
rect 10611 28228 10617 28230
rect 10588 28225 10617 28228
rect 11185 28224 11188 28230
rect 11214 28224 11217 28250
rect 12888 28245 12917 28248
rect 12888 28228 12894 28245
rect 12911 28244 12917 28245
rect 13071 28244 13074 28250
rect 12911 28230 13074 28244
rect 12911 28228 12917 28230
rect 12888 28225 12917 28228
rect 13071 28224 13074 28230
rect 13100 28224 13103 28250
rect 14497 28224 14500 28250
rect 14526 28244 14529 28250
rect 14636 28245 14665 28248
rect 14636 28244 14642 28245
rect 14526 28230 14642 28244
rect 14526 28224 14529 28230
rect 14636 28228 14642 28230
rect 14659 28228 14665 28245
rect 14636 28225 14665 28228
rect 15279 28224 15282 28250
rect 15308 28244 15311 28250
rect 15464 28245 15493 28248
rect 15464 28244 15470 28245
rect 15308 28230 15470 28244
rect 15308 28224 15311 28230
rect 15464 28228 15470 28230
rect 15487 28228 15493 28245
rect 15464 28225 15493 28228
rect 17303 28224 17306 28250
rect 17332 28244 17335 28250
rect 17350 28245 17379 28248
rect 17350 28244 17356 28245
rect 17332 28230 17356 28244
rect 17332 28224 17335 28230
rect 17350 28228 17356 28230
rect 17373 28228 17379 28245
rect 17350 28225 17379 28228
rect 17579 28224 17582 28250
rect 17608 28244 17611 28250
rect 17764 28245 17793 28248
rect 17764 28244 17770 28245
rect 17608 28230 17770 28244
rect 17608 28224 17611 28230
rect 17764 28228 17770 28230
rect 17787 28228 17793 28245
rect 17764 28225 17793 28228
rect 19373 28224 19376 28250
rect 19402 28224 19405 28250
rect 21075 28224 21078 28250
rect 21104 28224 21107 28250
rect 9299 28190 9302 28216
rect 9328 28210 9331 28216
rect 9760 28211 9789 28214
rect 9760 28210 9766 28211
rect 9328 28196 9766 28210
rect 9328 28190 9331 28196
rect 9760 28194 9766 28196
rect 9783 28210 9789 28211
rect 10220 28211 10249 28214
rect 10220 28210 10226 28211
rect 9783 28196 10226 28210
rect 9783 28194 9789 28196
rect 9760 28191 9789 28194
rect 10220 28194 10226 28196
rect 10243 28194 10249 28211
rect 11783 28210 11786 28216
rect 10220 28191 10249 28194
rect 10550 28196 11786 28210
rect 5436 28177 5465 28180
rect 5436 28160 5442 28177
rect 5459 28176 5465 28177
rect 5573 28176 5576 28182
rect 5459 28162 5576 28176
rect 5459 28160 5465 28162
rect 5436 28157 5465 28160
rect 5573 28156 5576 28162
rect 5602 28156 5605 28182
rect 8747 28156 8750 28182
rect 8776 28176 8779 28182
rect 8794 28177 8823 28180
rect 8794 28176 8800 28177
rect 8776 28162 8800 28176
rect 8776 28156 8779 28162
rect 8794 28160 8800 28162
rect 8817 28160 8823 28177
rect 8794 28157 8823 28160
rect 5481 28122 5484 28148
rect 5510 28122 5513 28148
rect 8802 28142 8816 28157
rect 8931 28156 8934 28182
rect 8960 28156 8963 28182
rect 9024 28177 9053 28180
rect 9024 28160 9030 28177
rect 9047 28176 9053 28177
rect 9115 28176 9118 28182
rect 9047 28162 9118 28176
rect 9047 28160 9053 28162
rect 9024 28157 9053 28160
rect 9115 28156 9118 28162
rect 9144 28156 9147 28182
rect 9668 28177 9697 28180
rect 9668 28160 9674 28177
rect 9691 28160 9697 28177
rect 9668 28157 9697 28160
rect 10128 28177 10157 28180
rect 10128 28160 10134 28177
rect 10151 28176 10157 28177
rect 10173 28176 10176 28182
rect 10151 28162 10176 28176
rect 10151 28160 10157 28162
rect 10128 28157 10157 28160
rect 9676 28142 9690 28157
rect 10173 28156 10176 28162
rect 10202 28156 10205 28182
rect 10266 28177 10295 28180
rect 10266 28160 10272 28177
rect 10289 28176 10295 28177
rect 10357 28176 10360 28182
rect 10289 28162 10360 28176
rect 10289 28160 10295 28162
rect 10266 28157 10295 28160
rect 10357 28156 10360 28162
rect 10386 28156 10389 28182
rect 10495 28156 10498 28182
rect 10524 28180 10527 28182
rect 10524 28177 10533 28180
rect 10527 28176 10533 28177
rect 10550 28176 10564 28196
rect 11783 28190 11786 28196
rect 11812 28190 11815 28216
rect 11968 28211 11997 28214
rect 11968 28194 11974 28211
rect 11991 28210 11997 28211
rect 12243 28210 12246 28216
rect 11991 28196 12246 28210
rect 11991 28194 11997 28196
rect 11968 28191 11997 28194
rect 12243 28190 12246 28196
rect 12272 28210 12275 28216
rect 15969 28210 15972 28216
rect 12272 28196 12910 28210
rect 12272 28190 12275 28196
rect 10527 28162 10564 28176
rect 10527 28160 10533 28162
rect 10524 28157 10533 28160
rect 10524 28156 10527 28157
rect 11001 28156 11004 28182
rect 11030 28176 11033 28182
rect 11830 28177 11859 28180
rect 11830 28176 11836 28177
rect 11030 28162 11836 28176
rect 11030 28156 11033 28162
rect 11830 28160 11836 28162
rect 11853 28160 11859 28177
rect 11830 28157 11859 28160
rect 12014 28177 12043 28180
rect 12014 28160 12020 28177
rect 12037 28176 12043 28177
rect 12381 28176 12384 28182
rect 12037 28162 12384 28176
rect 12037 28160 12043 28162
rect 12014 28157 12043 28160
rect 12381 28156 12384 28162
rect 12410 28156 12413 28182
rect 12896 28180 12910 28196
rect 13402 28196 14474 28210
rect 12796 28177 12825 28180
rect 12796 28160 12802 28177
rect 12819 28160 12825 28177
rect 12796 28157 12825 28160
rect 12888 28177 12917 28180
rect 12888 28160 12894 28177
rect 12911 28160 12917 28177
rect 12888 28157 12917 28160
rect 10680 28143 10709 28146
rect 10680 28142 10686 28143
rect 8802 28128 10686 28142
rect 10680 28126 10686 28128
rect 10703 28142 10709 28143
rect 10863 28142 10866 28148
rect 10703 28128 10866 28142
rect 10703 28126 10709 28128
rect 10680 28123 10709 28126
rect 10863 28122 10866 28128
rect 10892 28142 10895 28148
rect 11691 28142 11694 28148
rect 10892 28128 11694 28142
rect 10892 28122 10895 28128
rect 11691 28122 11694 28128
rect 11720 28142 11723 28148
rect 11738 28143 11767 28146
rect 11738 28142 11744 28143
rect 11720 28128 11744 28142
rect 11720 28122 11723 28128
rect 11738 28126 11744 28128
rect 11761 28126 11767 28143
rect 12804 28142 12818 28157
rect 13301 28156 13304 28182
rect 13330 28156 13333 28182
rect 13402 28180 13416 28196
rect 14460 28182 14474 28196
rect 15656 28196 15972 28210
rect 13394 28177 13423 28180
rect 13394 28160 13400 28177
rect 13417 28160 13423 28177
rect 13394 28157 13423 28160
rect 14313 28156 14316 28182
rect 14342 28156 14345 28182
rect 14359 28156 14362 28182
rect 14388 28176 14391 28182
rect 14388 28162 14410 28176
rect 14388 28156 14391 28162
rect 14451 28156 14454 28182
rect 14480 28156 14483 28182
rect 14497 28156 14500 28182
rect 14526 28156 14529 28182
rect 14543 28156 14546 28182
rect 14572 28180 14575 28182
rect 14572 28176 14576 28180
rect 14572 28162 14594 28176
rect 14572 28157 14576 28162
rect 14572 28156 14575 28157
rect 15463 28156 15466 28182
rect 15492 28156 15495 28182
rect 15656 28180 15670 28196
rect 15969 28190 15972 28196
rect 15998 28190 16001 28216
rect 17395 28190 17398 28216
rect 17424 28210 17427 28216
rect 18132 28211 18161 28214
rect 18132 28210 18138 28211
rect 17424 28196 18138 28210
rect 17424 28190 17427 28196
rect 18132 28194 18138 28196
rect 18155 28194 18161 28211
rect 18132 28191 18161 28194
rect 20707 28190 20710 28216
rect 20736 28190 20739 28216
rect 20845 28190 20848 28216
rect 20874 28190 20877 28216
rect 15648 28177 15677 28180
rect 15648 28160 15654 28177
rect 15671 28160 15677 28177
rect 15648 28157 15677 28160
rect 15831 28156 15834 28182
rect 15860 28156 15863 28182
rect 16705 28156 16708 28182
rect 16734 28176 16737 28182
rect 17073 28176 17076 28182
rect 16734 28162 17076 28176
rect 16734 28156 16737 28162
rect 17073 28156 17076 28162
rect 17102 28156 17105 28182
rect 17165 28156 17168 28182
rect 17194 28176 17197 28182
rect 17212 28177 17241 28180
rect 17212 28176 17218 28177
rect 17194 28162 17218 28176
rect 17194 28156 17197 28162
rect 17212 28160 17218 28162
rect 17235 28160 17241 28177
rect 17212 28157 17241 28160
rect 17257 28156 17260 28182
rect 17286 28176 17289 28182
rect 17856 28177 17885 28180
rect 17856 28176 17862 28177
rect 17286 28162 17862 28176
rect 17286 28156 17289 28162
rect 17856 28160 17862 28162
rect 17879 28160 17885 28177
rect 17856 28157 17885 28160
rect 18085 28156 18088 28182
rect 18114 28156 18117 28182
rect 18178 28177 18207 28180
rect 18178 28160 18184 28177
rect 18201 28160 18207 28177
rect 18178 28157 18207 28160
rect 18818 28177 18847 28180
rect 18818 28160 18824 28177
rect 18841 28176 18847 28177
rect 19005 28176 19008 28182
rect 18841 28162 19008 28176
rect 18841 28160 18847 28162
rect 18818 28157 18847 28160
rect 13348 28143 13377 28146
rect 13348 28142 13354 28143
rect 12804 28128 13354 28142
rect 11738 28123 11767 28126
rect 13348 28126 13354 28128
rect 13371 28126 13377 28143
rect 13348 28123 13377 28126
rect 14129 28122 14132 28148
rect 14158 28142 14161 28148
rect 14368 28142 14382 28156
rect 14158 28128 14382 28142
rect 17304 28143 17333 28146
rect 14158 28122 14161 28128
rect 17304 28126 17310 28143
rect 17327 28142 17333 28143
rect 17327 28128 17740 28142
rect 17327 28126 17333 28128
rect 17304 28123 17333 28126
rect 10127 28088 10130 28114
rect 10156 28088 10159 28114
rect 17441 28088 17444 28114
rect 17470 28108 17473 28114
rect 17672 28109 17701 28112
rect 17672 28108 17678 28109
rect 17470 28094 17678 28108
rect 17470 28088 17473 28094
rect 17672 28092 17678 28094
rect 17695 28092 17701 28109
rect 17726 28108 17740 28128
rect 17809 28122 17812 28148
rect 17838 28122 17841 28148
rect 17901 28122 17904 28148
rect 17930 28142 17933 28148
rect 18186 28142 18200 28157
rect 19005 28156 19008 28162
rect 19034 28156 19037 28182
rect 17930 28128 18200 28142
rect 17930 28122 17933 28128
rect 18683 28122 18686 28148
rect 18712 28122 18715 28148
rect 20155 28122 20158 28148
rect 20184 28142 20187 28148
rect 20202 28143 20231 28146
rect 20202 28142 20208 28143
rect 20184 28128 20208 28142
rect 20184 28122 20187 28128
rect 20202 28126 20208 28128
rect 20225 28126 20231 28143
rect 20202 28123 20231 28126
rect 20339 28122 20342 28148
rect 20368 28122 20371 28148
rect 18085 28108 18088 28114
rect 17726 28094 18088 28108
rect 17672 28089 17701 28092
rect 8655 28054 8658 28080
rect 8684 28074 8687 28080
rect 8863 28075 8892 28078
rect 8863 28074 8869 28075
rect 8684 28060 8869 28074
rect 8684 28054 8687 28060
rect 8863 28058 8869 28060
rect 8886 28058 8892 28075
rect 8863 28055 8892 28058
rect 10495 28054 10498 28080
rect 10524 28074 10527 28080
rect 10542 28075 10571 28078
rect 10542 28074 10548 28075
rect 10524 28060 10548 28074
rect 10524 28054 10527 28060
rect 10542 28058 10548 28060
rect 10565 28058 10571 28075
rect 17680 28074 17694 28089
rect 18085 28088 18088 28094
rect 18114 28088 18117 28114
rect 19235 28074 19238 28080
rect 17680 28060 19238 28074
rect 10542 28055 10571 28058
rect 19235 28054 19238 28060
rect 19264 28054 19267 28080
rect 3036 27992 29992 28040
rect 10173 27952 10176 27978
rect 10202 27972 10205 27978
rect 10450 27973 10479 27976
rect 10450 27972 10456 27973
rect 10202 27958 10456 27972
rect 10202 27952 10205 27958
rect 10450 27956 10456 27958
rect 10473 27956 10479 27973
rect 10450 27953 10479 27956
rect 17718 27973 17747 27976
rect 17718 27956 17724 27973
rect 17741 27972 17747 27973
rect 17809 27972 17812 27978
rect 17741 27958 17812 27972
rect 17741 27956 17747 27958
rect 17718 27953 17747 27956
rect 17809 27952 17812 27958
rect 17838 27952 17841 27978
rect 20339 27952 20342 27978
rect 20368 27952 20371 27978
rect 14451 27918 14454 27944
rect 14480 27938 14483 27944
rect 17396 27939 17425 27942
rect 17396 27938 17402 27939
rect 14480 27924 17402 27938
rect 14480 27918 14483 27924
rect 17396 27922 17402 27924
rect 17419 27922 17425 27939
rect 17396 27919 17425 27922
rect 17166 27905 17195 27908
rect 17166 27888 17172 27905
rect 17189 27904 17195 27905
rect 17211 27904 17214 27910
rect 17189 27890 17214 27904
rect 17189 27888 17195 27890
rect 17166 27885 17195 27888
rect 17211 27884 17214 27890
rect 17240 27884 17243 27910
rect 17441 27884 17444 27910
rect 17470 27884 17473 27910
rect 20615 27884 20618 27910
rect 20644 27884 20647 27910
rect 10403 27850 10406 27876
rect 10432 27850 10435 27876
rect 10495 27850 10498 27876
rect 10524 27850 10527 27876
rect 11600 27871 11629 27874
rect 11600 27854 11606 27871
rect 11623 27870 11629 27871
rect 11645 27870 11648 27876
rect 11623 27856 11648 27870
rect 11623 27854 11629 27856
rect 11600 27851 11629 27854
rect 11645 27850 11648 27856
rect 11674 27850 11677 27876
rect 11692 27871 11721 27874
rect 11692 27854 11698 27871
rect 11715 27870 11721 27871
rect 11783 27870 11786 27876
rect 11715 27856 11786 27870
rect 11715 27854 11721 27856
rect 11692 27851 11721 27854
rect 11783 27850 11786 27856
rect 11812 27870 11815 27876
rect 12060 27871 12089 27874
rect 11812 27856 11990 27870
rect 11812 27850 11815 27856
rect 11599 27782 11602 27808
rect 11628 27802 11631 27808
rect 11976 27806 11990 27856
rect 12060 27854 12066 27871
rect 12083 27870 12089 27871
rect 12105 27870 12108 27876
rect 12083 27856 12108 27870
rect 12083 27854 12089 27856
rect 12060 27851 12089 27854
rect 12105 27850 12108 27856
rect 12134 27850 12137 27876
rect 12381 27850 12384 27876
rect 12410 27870 12413 27876
rect 14497 27870 14500 27876
rect 12410 27856 14500 27870
rect 12410 27850 12413 27856
rect 14497 27850 14500 27856
rect 14526 27870 14529 27876
rect 15279 27870 15282 27876
rect 14526 27856 15282 27870
rect 14526 27850 14529 27856
rect 15279 27850 15282 27856
rect 15308 27850 15311 27876
rect 17258 27871 17287 27874
rect 17258 27854 17264 27871
rect 17281 27854 17287 27871
rect 17258 27851 17287 27854
rect 17266 27836 17280 27851
rect 17671 27850 17674 27876
rect 17700 27850 17703 27876
rect 17764 27871 17793 27874
rect 17764 27854 17770 27871
rect 17787 27870 17793 27871
rect 18085 27870 18088 27876
rect 17787 27856 18088 27870
rect 17787 27854 17793 27856
rect 17764 27851 17793 27854
rect 18085 27850 18088 27856
rect 18114 27850 18117 27876
rect 18683 27850 18686 27876
rect 18712 27870 18715 27876
rect 19097 27870 19100 27876
rect 18712 27856 19100 27870
rect 18712 27850 18715 27856
rect 19097 27850 19100 27856
rect 19126 27850 19129 27876
rect 19622 27871 19651 27874
rect 19622 27870 19628 27871
rect 19382 27856 19628 27870
rect 17718 27837 17747 27840
rect 17718 27836 17724 27837
rect 17266 27822 17724 27836
rect 17718 27820 17724 27822
rect 17741 27820 17747 27837
rect 17718 27817 17747 27820
rect 18729 27816 18732 27842
rect 18758 27836 18761 27842
rect 18807 27837 18836 27840
rect 18807 27836 18813 27837
rect 18758 27822 18813 27836
rect 18758 27816 18761 27822
rect 18807 27820 18813 27822
rect 18830 27820 18836 27837
rect 18807 27817 18836 27820
rect 11646 27803 11675 27806
rect 11646 27802 11652 27803
rect 11628 27788 11652 27802
rect 11628 27782 11631 27788
rect 11646 27786 11652 27788
rect 11669 27786 11675 27803
rect 11646 27783 11675 27786
rect 11968 27803 11997 27806
rect 11968 27786 11974 27803
rect 11991 27786 11997 27803
rect 11968 27783 11997 27786
rect 17441 27782 17444 27808
rect 17470 27802 17473 27808
rect 17901 27802 17904 27808
rect 17470 27788 17904 27802
rect 17470 27782 17473 27788
rect 17901 27782 17904 27788
rect 17930 27782 17933 27808
rect 19005 27782 19008 27808
rect 19034 27802 19037 27808
rect 19382 27806 19396 27856
rect 19622 27854 19628 27856
rect 19645 27854 19651 27871
rect 19622 27851 19651 27854
rect 20524 27871 20553 27874
rect 20524 27854 20530 27871
rect 20547 27870 20553 27871
rect 21075 27870 21078 27876
rect 20547 27856 21078 27870
rect 20547 27854 20553 27856
rect 20524 27851 20553 27854
rect 21075 27850 21078 27856
rect 21104 27850 21107 27876
rect 19374 27803 19403 27806
rect 19374 27802 19380 27803
rect 19034 27788 19380 27802
rect 19034 27782 19037 27788
rect 19374 27786 19380 27788
rect 19397 27786 19403 27803
rect 19374 27783 19403 27786
rect 19465 27782 19468 27808
rect 19494 27802 19497 27808
rect 19673 27803 19702 27806
rect 19673 27802 19679 27803
rect 19494 27788 19679 27802
rect 19494 27782 19497 27788
rect 19673 27786 19679 27788
rect 19696 27786 19702 27803
rect 19673 27783 19702 27786
rect 20569 27782 20572 27808
rect 20598 27782 20601 27808
rect 3036 27720 29992 27768
rect 6769 27680 6772 27706
rect 6798 27680 6801 27706
rect 12105 27680 12108 27706
rect 12134 27700 12137 27706
rect 12134 27686 14612 27700
rect 12134 27680 12137 27686
rect 4727 27667 4756 27670
rect 4727 27650 4733 27667
rect 4750 27666 4756 27667
rect 4791 27666 4794 27672
rect 4750 27652 4794 27666
rect 4750 27650 4756 27652
rect 4727 27647 4756 27650
rect 4791 27646 4794 27652
rect 4820 27646 4823 27672
rect 6778 27666 6792 27680
rect 6456 27652 6792 27666
rect 4677 27633 4706 27636
rect 4677 27616 4683 27633
rect 4700 27632 4706 27633
rect 5067 27632 5070 27638
rect 4700 27618 5070 27632
rect 4700 27616 4706 27618
rect 4677 27613 4706 27616
rect 5067 27612 5070 27618
rect 5096 27612 5099 27638
rect 6456 27636 6470 27652
rect 6953 27646 6956 27672
rect 6982 27646 6985 27672
rect 7367 27646 7370 27672
rect 7396 27646 7399 27672
rect 8655 27646 8658 27672
rect 8684 27666 8687 27672
rect 10541 27666 10544 27672
rect 8684 27652 10544 27666
rect 8684 27646 8687 27652
rect 6448 27633 6477 27636
rect 6448 27616 6454 27633
rect 6471 27616 6477 27633
rect 6448 27613 6477 27616
rect 6540 27633 6569 27636
rect 6540 27616 6546 27633
rect 6563 27632 6569 27633
rect 6677 27632 6680 27638
rect 6563 27618 6680 27632
rect 6563 27616 6569 27618
rect 6540 27613 6569 27616
rect 6677 27612 6680 27618
rect 6706 27612 6709 27638
rect 6770 27633 6799 27636
rect 6770 27616 6776 27633
rect 6793 27632 6799 27633
rect 6962 27632 6976 27646
rect 7183 27632 7186 27638
rect 6793 27618 7186 27632
rect 6793 27616 6799 27618
rect 6770 27613 6799 27616
rect 7183 27612 7186 27618
rect 7212 27612 7215 27638
rect 7284 27618 7666 27632
rect 4515 27578 4518 27604
rect 4544 27578 4547 27604
rect 5527 27578 5530 27604
rect 5556 27602 5559 27604
rect 5556 27599 5580 27602
rect 5556 27582 5557 27599
rect 5574 27582 5580 27599
rect 5556 27579 5580 27582
rect 6908 27599 6937 27602
rect 6908 27582 6914 27599
rect 6931 27598 6937 27599
rect 6953 27598 6956 27604
rect 6931 27584 6956 27598
rect 6931 27582 6937 27584
rect 6908 27579 6937 27582
rect 5556 27578 5559 27579
rect 6953 27578 6956 27584
rect 6982 27578 6985 27604
rect 7284 27598 7298 27618
rect 7146 27584 7298 27598
rect 7322 27599 7351 27602
rect 6816 27565 6845 27568
rect 6816 27548 6822 27565
rect 6839 27564 6845 27565
rect 7146 27564 7160 27584
rect 7322 27582 7328 27599
rect 7345 27598 7351 27599
rect 7597 27598 7600 27604
rect 7345 27584 7600 27598
rect 7345 27582 7351 27584
rect 7322 27579 7351 27582
rect 7597 27578 7600 27584
rect 7626 27578 7629 27604
rect 7652 27598 7666 27618
rect 10265 27612 10268 27638
rect 10294 27612 10297 27638
rect 10412 27636 10426 27652
rect 10541 27646 10544 27652
rect 10570 27646 10573 27672
rect 11645 27646 11648 27672
rect 11674 27666 11677 27672
rect 14543 27666 14546 27672
rect 11674 27652 14546 27666
rect 11674 27646 11677 27652
rect 14543 27646 14546 27652
rect 14572 27646 14575 27672
rect 10404 27633 10433 27636
rect 10404 27616 10410 27633
rect 10427 27616 10433 27633
rect 10404 27613 10433 27616
rect 10450 27633 10479 27636
rect 10450 27616 10456 27633
rect 10473 27632 10479 27633
rect 11001 27632 11004 27638
rect 10473 27618 11004 27632
rect 10473 27616 10479 27618
rect 10450 27613 10479 27616
rect 11001 27612 11004 27618
rect 11030 27632 11033 27638
rect 11600 27633 11629 27636
rect 11600 27632 11606 27633
rect 11030 27618 11606 27632
rect 11030 27612 11033 27618
rect 11600 27616 11606 27618
rect 11623 27616 11629 27633
rect 11600 27613 11629 27616
rect 11691 27612 11694 27638
rect 11720 27612 11723 27638
rect 11921 27612 11924 27638
rect 11950 27632 11953 27638
rect 11968 27633 11997 27636
rect 11968 27632 11974 27633
rect 11950 27618 11974 27632
rect 11950 27612 11953 27618
rect 11968 27616 11974 27618
rect 11991 27616 11997 27633
rect 11968 27613 11997 27616
rect 12105 27612 12108 27638
rect 12134 27612 12137 27638
rect 12243 27612 12246 27638
rect 12272 27612 12275 27638
rect 13347 27612 13350 27638
rect 13376 27612 13379 27638
rect 13393 27612 13396 27638
rect 13422 27632 13425 27638
rect 13440 27633 13469 27636
rect 13440 27632 13446 27633
rect 13422 27618 13446 27632
rect 13422 27612 13425 27618
rect 13440 27616 13446 27618
rect 13463 27616 13469 27633
rect 13440 27613 13469 27616
rect 13486 27633 13515 27636
rect 13486 27616 13492 27633
rect 13509 27632 13515 27633
rect 13577 27632 13580 27638
rect 13509 27618 13580 27632
rect 13509 27616 13515 27618
rect 13486 27613 13515 27616
rect 13577 27612 13580 27618
rect 13606 27612 13609 27638
rect 14598 27632 14612 27686
rect 15877 27646 15880 27672
rect 15906 27646 15909 27672
rect 17671 27646 17674 27672
rect 17700 27666 17703 27672
rect 18408 27667 18437 27670
rect 18408 27666 18414 27667
rect 17700 27652 18414 27666
rect 17700 27646 17703 27652
rect 15141 27632 15144 27638
rect 14598 27618 15144 27632
rect 15141 27612 15144 27618
rect 15170 27612 15173 27638
rect 15279 27612 15282 27638
rect 15308 27612 15311 27638
rect 15694 27633 15723 27636
rect 15694 27616 15700 27633
rect 15717 27632 15723 27633
rect 15739 27632 15742 27638
rect 15717 27618 15742 27632
rect 15717 27616 15723 27618
rect 15694 27613 15723 27616
rect 15739 27612 15742 27618
rect 15768 27612 15771 27638
rect 15786 27633 15815 27636
rect 15786 27616 15792 27633
rect 15809 27632 15815 27633
rect 15886 27632 15900 27646
rect 15809 27618 15900 27632
rect 15809 27616 15815 27618
rect 15786 27613 15815 27616
rect 17993 27612 17996 27638
rect 18022 27612 18025 27638
rect 18094 27636 18108 27652
rect 18408 27650 18414 27652
rect 18431 27650 18437 27667
rect 18408 27647 18437 27650
rect 18914 27667 18943 27670
rect 18914 27650 18920 27667
rect 18937 27666 18943 27667
rect 19235 27666 19238 27672
rect 18937 27652 19238 27666
rect 18937 27650 18943 27652
rect 18914 27647 18943 27650
rect 19235 27646 19238 27652
rect 19264 27646 19267 27672
rect 18086 27633 18115 27636
rect 18086 27616 18092 27633
rect 18109 27616 18115 27633
rect 18453 27632 18456 27638
rect 18443 27618 18456 27632
rect 18086 27613 18115 27616
rect 18453 27612 18456 27618
rect 18482 27612 18485 27638
rect 19005 27612 19008 27638
rect 19034 27612 19037 27638
rect 7689 27598 7692 27604
rect 7652 27584 7692 27598
rect 7689 27578 7692 27584
rect 7718 27578 7721 27604
rect 12335 27578 12338 27604
rect 12364 27578 12367 27604
rect 15372 27599 15401 27602
rect 15372 27582 15378 27599
rect 15395 27582 15401 27599
rect 15372 27579 15401 27582
rect 6839 27550 7160 27564
rect 7184 27565 7213 27568
rect 6839 27548 6845 27550
rect 6816 27545 6845 27548
rect 7184 27548 7190 27565
rect 7207 27564 7213 27565
rect 7735 27564 7738 27570
rect 7207 27550 7738 27564
rect 7207 27548 7213 27550
rect 7184 27545 7213 27548
rect 7735 27544 7738 27550
rect 7764 27544 7767 27570
rect 10403 27544 10406 27570
rect 10432 27564 10435 27570
rect 10633 27564 10636 27570
rect 10432 27550 10636 27564
rect 10432 27544 10435 27550
rect 10633 27544 10636 27550
rect 10662 27564 10665 27570
rect 13301 27564 13304 27570
rect 10662 27550 13304 27564
rect 10662 27544 10665 27550
rect 13301 27544 13304 27550
rect 13330 27544 13333 27570
rect 15380 27564 15394 27579
rect 15463 27578 15466 27604
rect 15492 27578 15495 27604
rect 18462 27598 18476 27612
rect 19098 27599 19127 27602
rect 19098 27598 19104 27599
rect 18462 27584 19104 27598
rect 19098 27582 19104 27584
rect 19121 27582 19127 27599
rect 19098 27579 19127 27582
rect 15740 27565 15769 27568
rect 15740 27564 15746 27565
rect 15380 27550 15746 27564
rect 15740 27548 15746 27550
rect 15763 27548 15769 27565
rect 15740 27545 15769 27548
rect 18085 27544 18088 27570
rect 18114 27564 18117 27570
rect 18316 27565 18345 27568
rect 18316 27564 18322 27565
rect 18114 27550 18322 27564
rect 18114 27544 18117 27550
rect 18316 27548 18322 27550
rect 18339 27564 18345 27565
rect 18361 27564 18364 27570
rect 18339 27550 18364 27564
rect 18339 27548 18345 27550
rect 18316 27545 18345 27548
rect 18361 27544 18364 27550
rect 18390 27544 18393 27570
rect 18775 27564 18778 27570
rect 18508 27550 18778 27564
rect 6355 27510 6358 27536
rect 6384 27530 6387 27536
rect 6494 27531 6523 27534
rect 6494 27530 6500 27531
rect 6384 27516 6500 27530
rect 6384 27510 6387 27516
rect 6494 27514 6500 27516
rect 6517 27514 6523 27531
rect 6494 27511 6523 27514
rect 7230 27531 7259 27534
rect 7230 27514 7236 27531
rect 7253 27530 7259 27531
rect 7643 27530 7646 27536
rect 7253 27516 7646 27530
rect 7253 27514 7259 27516
rect 7230 27511 7259 27514
rect 7643 27510 7646 27516
rect 7672 27510 7675 27536
rect 13255 27510 13258 27536
rect 13284 27530 13287 27536
rect 13348 27531 13377 27534
rect 13348 27530 13354 27531
rect 13284 27516 13354 27530
rect 13284 27510 13287 27516
rect 13348 27514 13354 27516
rect 13371 27514 13377 27531
rect 13348 27511 13377 27514
rect 18040 27531 18069 27534
rect 18040 27514 18046 27531
rect 18063 27530 18069 27531
rect 18508 27530 18522 27550
rect 18775 27544 18778 27550
rect 18804 27544 18807 27570
rect 18063 27516 18522 27530
rect 18546 27531 18575 27534
rect 18063 27514 18069 27516
rect 18040 27511 18069 27514
rect 18546 27514 18552 27531
rect 18569 27530 18575 27531
rect 19373 27530 19376 27536
rect 18569 27516 19376 27530
rect 18569 27514 18575 27516
rect 18546 27511 18575 27514
rect 19373 27510 19376 27516
rect 19402 27510 19405 27536
rect 3036 27448 29992 27496
rect 6723 27428 6726 27434
rect 5352 27414 6726 27428
rect 4515 27306 4518 27332
rect 4544 27326 4547 27332
rect 4699 27326 4702 27332
rect 4544 27312 4702 27326
rect 4544 27306 4547 27312
rect 4699 27306 4702 27312
rect 4728 27326 4731 27332
rect 5352 27330 5366 27414
rect 6723 27408 6726 27414
rect 6752 27408 6755 27434
rect 18729 27408 18732 27434
rect 18758 27408 18761 27434
rect 19465 27428 19468 27434
rect 19152 27414 19468 27428
rect 6953 27374 6956 27400
rect 6982 27394 6985 27400
rect 8747 27394 8750 27400
rect 6982 27380 8750 27394
rect 6982 27374 6985 27380
rect 8747 27374 8750 27380
rect 8776 27374 8779 27400
rect 14957 27374 14960 27400
rect 14986 27374 14989 27400
rect 19152 27394 19166 27414
rect 19465 27408 19468 27414
rect 19494 27408 19497 27434
rect 20179 27429 20208 27432
rect 20179 27412 20185 27429
rect 20202 27428 20208 27429
rect 20569 27428 20572 27434
rect 20202 27414 20572 27428
rect 20202 27412 20208 27414
rect 20179 27409 20208 27412
rect 20569 27408 20572 27414
rect 20598 27408 20601 27434
rect 18646 27380 19166 27394
rect 6263 27340 6266 27366
rect 6292 27360 6295 27366
rect 6379 27361 6408 27364
rect 6379 27360 6385 27361
rect 6292 27346 6385 27360
rect 6292 27340 6295 27346
rect 6379 27344 6385 27346
rect 6402 27344 6408 27361
rect 6379 27341 6408 27344
rect 7367 27340 7370 27366
rect 7396 27360 7399 27366
rect 7552 27361 7581 27364
rect 7552 27360 7558 27361
rect 7396 27346 7558 27360
rect 7396 27340 7399 27346
rect 7552 27344 7558 27346
rect 7575 27344 7581 27361
rect 7552 27341 7581 27344
rect 7643 27340 7646 27366
rect 7672 27340 7675 27366
rect 5344 27327 5373 27330
rect 5344 27326 5350 27327
rect 4728 27312 5350 27326
rect 4728 27306 4731 27312
rect 5344 27310 5350 27312
rect 5367 27310 5373 27327
rect 5344 27307 5373 27310
rect 5505 27327 5534 27330
rect 5505 27310 5511 27327
rect 5528 27326 5534 27327
rect 6033 27326 6036 27332
rect 5528 27312 6036 27326
rect 5528 27310 5534 27312
rect 5505 27307 5534 27310
rect 6033 27306 6036 27312
rect 6062 27306 6065 27332
rect 7505 27306 7508 27332
rect 7534 27306 7537 27332
rect 7597 27306 7600 27332
rect 7626 27326 7629 27332
rect 7626 27312 8172 27326
rect 7626 27306 7629 27312
rect 5555 27293 5584 27296
rect 5555 27276 5561 27293
rect 5578 27292 5584 27293
rect 5619 27292 5622 27298
rect 5578 27278 5622 27292
rect 5578 27276 5584 27278
rect 5555 27273 5584 27276
rect 5619 27272 5622 27278
rect 5648 27272 5651 27298
rect 8158 27264 8172 27312
rect 8655 27306 8658 27332
rect 8684 27306 8687 27332
rect 8756 27326 8770 27374
rect 9530 27361 9559 27364
rect 9530 27344 9536 27361
rect 9553 27360 9559 27361
rect 10265 27360 10268 27366
rect 9553 27346 10268 27360
rect 9553 27344 9559 27346
rect 9530 27341 9559 27344
rect 10265 27340 10268 27346
rect 10294 27340 10297 27366
rect 8794 27327 8823 27330
rect 8794 27326 8800 27327
rect 8756 27312 8800 27326
rect 8794 27310 8800 27312
rect 8817 27310 8823 27327
rect 8794 27307 8823 27310
rect 9345 27306 9348 27332
rect 9374 27306 9377 27332
rect 9713 27306 9716 27332
rect 9742 27306 9745 27332
rect 13117 27306 13120 27332
rect 13146 27306 13149 27332
rect 13255 27330 13258 27332
rect 13252 27326 13258 27330
rect 13235 27312 13258 27326
rect 13252 27307 13258 27312
rect 13255 27306 13258 27307
rect 13284 27306 13287 27332
rect 15096 27327 15125 27330
rect 15096 27310 15102 27327
rect 15119 27326 15125 27327
rect 16429 27326 16432 27332
rect 15119 27312 16432 27326
rect 15119 27310 15125 27312
rect 15096 27307 15125 27310
rect 16429 27306 16432 27312
rect 16458 27306 16461 27332
rect 16476 27327 16505 27330
rect 16476 27310 16482 27327
rect 16499 27310 16505 27327
rect 16476 27307 16505 27310
rect 16568 27327 16597 27330
rect 16568 27310 16574 27327
rect 16591 27326 16597 27327
rect 17165 27326 17168 27332
rect 16591 27312 17168 27326
rect 16591 27310 16597 27312
rect 16568 27307 16597 27310
rect 8747 27272 8750 27298
rect 8776 27272 8779 27298
rect 14589 27272 14592 27298
rect 14618 27292 14621 27298
rect 14958 27293 14987 27296
rect 14958 27292 14964 27293
rect 14618 27278 14964 27292
rect 14618 27272 14621 27278
rect 14958 27276 14964 27278
rect 14981 27292 14987 27293
rect 16484 27292 16498 27307
rect 17165 27306 17168 27312
rect 17194 27306 17197 27332
rect 18646 27330 18660 27380
rect 18775 27340 18778 27366
rect 18804 27340 18807 27366
rect 18638 27327 18667 27330
rect 18638 27310 18644 27327
rect 18661 27310 18667 27327
rect 18638 27307 18667 27310
rect 18684 27327 18713 27330
rect 18684 27310 18690 27327
rect 18707 27310 18713 27327
rect 18684 27307 18713 27310
rect 14981 27278 15118 27292
rect 16484 27278 16590 27292
rect 14981 27276 14987 27278
rect 14958 27273 14987 27276
rect 15104 27264 15118 27278
rect 16576 27264 16590 27278
rect 6769 27238 6772 27264
rect 6798 27258 6801 27264
rect 7045 27258 7048 27264
rect 6798 27244 7048 27258
rect 6798 27238 6801 27244
rect 7045 27238 7048 27244
rect 7074 27238 7077 27264
rect 7413 27238 7416 27264
rect 7442 27238 7445 27264
rect 8149 27238 8152 27264
rect 8178 27258 8181 27264
rect 9300 27259 9329 27262
rect 9300 27258 9306 27259
rect 8178 27244 9306 27258
rect 8178 27238 8181 27244
rect 9300 27242 9306 27244
rect 9323 27242 9329 27259
rect 9300 27239 9329 27242
rect 13255 27238 13258 27264
rect 13284 27258 13287 27264
rect 13393 27258 13396 27264
rect 13284 27244 13396 27258
rect 13284 27238 13287 27244
rect 13393 27238 13396 27244
rect 13422 27258 13425 27264
rect 13808 27259 13837 27262
rect 13808 27258 13814 27259
rect 13422 27244 13814 27258
rect 13422 27238 13425 27244
rect 13808 27242 13814 27244
rect 13831 27242 13837 27259
rect 13808 27239 13837 27242
rect 15049 27238 15052 27264
rect 15078 27238 15081 27264
rect 15095 27238 15098 27264
rect 15124 27238 15127 27264
rect 16475 27238 16478 27264
rect 16504 27258 16507 27264
rect 16522 27259 16551 27262
rect 16522 27258 16528 27259
rect 16504 27244 16528 27258
rect 16504 27238 16507 27244
rect 16522 27242 16528 27244
rect 16545 27242 16551 27259
rect 16522 27239 16551 27242
rect 16567 27238 16570 27264
rect 16596 27258 16599 27264
rect 18692 27258 18706 27307
rect 19097 27306 19100 27332
rect 19126 27326 19129 27332
rect 19144 27327 19173 27330
rect 19144 27326 19150 27327
rect 19126 27312 19150 27326
rect 19126 27306 19129 27312
rect 19144 27310 19150 27312
rect 19167 27310 19173 27327
rect 19144 27307 19173 27310
rect 19305 27327 19334 27330
rect 19305 27310 19311 27327
rect 19328 27326 19334 27327
rect 19419 27326 19422 27332
rect 19328 27312 19422 27326
rect 19328 27310 19334 27312
rect 19305 27307 19334 27310
rect 19419 27306 19422 27312
rect 19448 27306 19451 27332
rect 19373 27296 19376 27298
rect 19355 27293 19376 27296
rect 19355 27276 19361 27293
rect 19355 27273 19376 27276
rect 19373 27272 19376 27273
rect 19402 27272 19405 27298
rect 16596 27244 18706 27258
rect 16596 27238 16599 27244
rect 3036 27176 29992 27224
rect 5573 27160 5576 27162
rect 5551 27157 5576 27160
rect 5551 27140 5557 27157
rect 5574 27140 5576 27157
rect 5551 27137 5576 27140
rect 5573 27136 5576 27137
rect 5602 27136 5605 27162
rect 6033 27136 6036 27162
rect 6062 27136 6065 27162
rect 6263 27136 6266 27162
rect 6292 27136 6295 27162
rect 7735 27136 7738 27162
rect 7764 27160 7767 27162
rect 7764 27157 7788 27160
rect 7764 27140 7765 27157
rect 7782 27140 7788 27157
rect 7764 27137 7788 27140
rect 7764 27136 7767 27137
rect 11921 27136 11924 27162
rect 11950 27136 11953 27162
rect 13347 27136 13350 27162
rect 13376 27156 13379 27162
rect 13486 27157 13515 27160
rect 13486 27156 13492 27157
rect 13376 27142 13492 27156
rect 13376 27136 13379 27142
rect 13486 27140 13492 27142
rect 13509 27140 13515 27157
rect 13486 27137 13515 27140
rect 15141 27136 15144 27162
rect 15170 27156 15173 27162
rect 15280 27157 15309 27160
rect 15280 27156 15286 27157
rect 15170 27142 15286 27156
rect 15170 27136 15173 27142
rect 15280 27140 15286 27142
rect 15303 27140 15309 27157
rect 15280 27137 15309 27140
rect 17993 27136 17996 27162
rect 18022 27156 18025 27162
rect 18362 27157 18391 27160
rect 18362 27156 18368 27157
rect 18022 27142 18368 27156
rect 18022 27136 18025 27142
rect 18362 27140 18368 27142
rect 18385 27140 18391 27157
rect 18362 27137 18391 27140
rect 5619 27102 5622 27128
rect 5648 27122 5651 27128
rect 6769 27122 6772 27128
rect 5648 27108 6772 27122
rect 5648 27102 5651 27108
rect 6769 27102 6772 27108
rect 6798 27122 6801 27128
rect 6931 27123 6960 27126
rect 6931 27122 6937 27123
rect 6798 27108 6937 27122
rect 6798 27102 6801 27108
rect 6931 27106 6937 27108
rect 6954 27106 6960 27123
rect 6931 27103 6960 27106
rect 8149 27102 8152 27128
rect 8178 27102 8181 27128
rect 8195 27102 8198 27128
rect 8224 27122 8227 27128
rect 9345 27122 9348 27128
rect 8224 27108 9348 27122
rect 8224 27102 8227 27108
rect 9345 27102 9348 27108
rect 9374 27122 9377 27128
rect 9392 27123 9421 27126
rect 9392 27122 9398 27123
rect 9374 27108 9398 27122
rect 9374 27102 9377 27108
rect 9392 27106 9398 27108
rect 9415 27106 9421 27123
rect 9392 27103 9421 27106
rect 10633 27102 10636 27128
rect 10662 27102 10665 27128
rect 10725 27102 10728 27128
rect 10754 27126 10757 27128
rect 10754 27123 10763 27126
rect 10757 27106 10763 27123
rect 12381 27122 12384 27128
rect 10754 27103 10763 27106
rect 11976 27108 12384 27122
rect 10754 27102 10757 27103
rect 4653 27068 4656 27094
rect 4682 27092 4685 27094
rect 4682 27089 4700 27092
rect 4694 27072 4700 27089
rect 4682 27069 4700 27072
rect 4715 27089 4744 27092
rect 4715 27072 4721 27089
rect 4738 27088 4744 27089
rect 4791 27088 4794 27094
rect 4738 27074 4794 27088
rect 4738 27072 4744 27074
rect 4715 27069 4744 27072
rect 4682 27068 4685 27069
rect 4791 27068 4794 27074
rect 4820 27088 4823 27094
rect 5251 27088 5254 27094
rect 4820 27074 5254 27088
rect 4820 27068 4823 27074
rect 5251 27068 5254 27074
rect 5280 27068 5283 27094
rect 6217 27068 6220 27094
rect 6246 27068 6249 27094
rect 6723 27068 6726 27094
rect 6752 27068 6755 27094
rect 6885 27089 6914 27092
rect 6885 27072 6891 27089
rect 6908 27088 6914 27089
rect 7413 27088 7416 27094
rect 6908 27074 7416 27088
rect 6908 27072 6914 27074
rect 6885 27069 6914 27072
rect 7413 27068 7416 27074
rect 7442 27068 7445 27094
rect 8242 27089 8271 27092
rect 8242 27072 8248 27089
rect 8265 27088 8271 27089
rect 8747 27088 8750 27094
rect 8265 27074 8750 27088
rect 8265 27072 8271 27074
rect 8242 27069 8271 27072
rect 8747 27068 8750 27074
rect 8776 27088 8779 27094
rect 8886 27089 8915 27092
rect 8886 27088 8892 27089
rect 8776 27074 8892 27088
rect 8776 27068 8779 27074
rect 8886 27072 8892 27074
rect 8909 27088 8915 27089
rect 9254 27089 9283 27092
rect 9254 27088 9260 27089
rect 8909 27074 9260 27088
rect 8909 27072 8915 27074
rect 8886 27069 8915 27072
rect 9254 27072 9260 27074
rect 9277 27072 9283 27089
rect 9254 27069 9283 27072
rect 11830 27089 11859 27092
rect 11830 27072 11836 27089
rect 11853 27088 11859 27089
rect 11921 27088 11924 27094
rect 11853 27074 11924 27088
rect 11853 27072 11859 27074
rect 11830 27069 11859 27072
rect 11921 27068 11924 27074
rect 11950 27068 11953 27094
rect 11976 27092 11990 27108
rect 12381 27102 12384 27108
rect 12410 27102 12413 27128
rect 14589 27122 14592 27128
rect 13103 27108 14592 27122
rect 11968 27089 11997 27092
rect 11968 27072 11974 27089
rect 11991 27072 11997 27089
rect 11968 27069 11997 27072
rect 12198 27089 12227 27092
rect 12198 27072 12204 27089
rect 12221 27072 12227 27089
rect 12198 27069 12227 27072
rect 4515 27034 4518 27060
rect 4544 27034 4547 27060
rect 6264 27055 6293 27058
rect 6264 27038 6270 27055
rect 6287 27038 6293 27055
rect 6264 27035 6293 27038
rect 6272 26986 6286 27035
rect 6355 27034 6358 27060
rect 6384 27034 6387 27060
rect 7597 27034 7600 27060
rect 7626 27054 7629 27060
rect 8932 27055 8961 27058
rect 8932 27054 8938 27055
rect 7626 27040 8938 27054
rect 7626 27034 7629 27040
rect 7413 26986 7416 26992
rect 6272 26972 7416 26986
rect 7413 26966 7416 26972
rect 7442 26966 7445 26992
rect 8333 26966 8336 26992
rect 8362 26966 8365 26992
rect 8655 26966 8658 26992
rect 8684 26986 8687 26992
rect 8794 26987 8823 26990
rect 8794 26986 8800 26987
rect 8684 26972 8800 26986
rect 8684 26966 8687 26972
rect 8794 26970 8800 26972
rect 8817 26970 8823 26987
rect 8894 26986 8908 27040
rect 8932 27038 8938 27040
rect 8955 27038 8961 27055
rect 8932 27035 8961 27038
rect 8978 27055 9007 27058
rect 8978 27038 8984 27055
rect 9001 27054 9007 27055
rect 9392 27055 9421 27058
rect 9392 27054 9398 27055
rect 9001 27040 9398 27054
rect 9001 27038 9007 27040
rect 8978 27035 9007 27038
rect 9392 27038 9398 27040
rect 9415 27038 9421 27055
rect 12206 27054 12220 27069
rect 12289 27068 12292 27094
rect 12318 27088 12321 27094
rect 13103 27088 13117 27108
rect 14589 27102 14592 27108
rect 14618 27102 14621 27128
rect 14724 27123 14753 27126
rect 14724 27106 14730 27123
rect 14747 27122 14753 27123
rect 14957 27122 14960 27128
rect 14747 27108 14960 27122
rect 14747 27106 14753 27108
rect 14724 27103 14753 27106
rect 14957 27102 14960 27108
rect 14986 27102 14989 27128
rect 15003 27102 15006 27128
rect 15032 27122 15035 27128
rect 15463 27122 15466 27128
rect 15032 27108 15466 27122
rect 15032 27102 15035 27108
rect 15463 27102 15466 27108
rect 15492 27122 15495 27128
rect 16384 27123 16413 27126
rect 16384 27122 16390 27123
rect 15492 27108 16390 27122
rect 15492 27102 15495 27108
rect 16384 27106 16390 27108
rect 16407 27122 16413 27123
rect 16567 27122 16570 27128
rect 16407 27108 16570 27122
rect 16407 27106 16413 27108
rect 16384 27103 16413 27106
rect 16567 27102 16570 27108
rect 16596 27102 16599 27128
rect 20707 27102 20710 27128
rect 20736 27102 20739 27128
rect 21305 27122 21308 27128
rect 21045 27108 21308 27122
rect 21305 27102 21308 27108
rect 21334 27102 21337 27128
rect 12318 27074 13117 27088
rect 12318 27068 12321 27074
rect 13301 27068 13304 27094
rect 13330 27088 13333 27094
rect 13330 27074 13508 27088
rect 13330 27068 13333 27074
rect 9392 27035 9421 27038
rect 11838 27040 12220 27054
rect 9300 27021 9329 27024
rect 9300 27004 9306 27021
rect 9323 27020 9329 27021
rect 9713 27020 9716 27026
rect 9323 27006 9716 27020
rect 9323 27004 9329 27006
rect 9300 27001 9329 27004
rect 9308 26986 9322 27001
rect 9713 27000 9716 27006
rect 9742 27000 9745 27026
rect 11599 27020 11602 27026
rect 10734 27006 11602 27020
rect 8894 26972 9322 26986
rect 8794 26967 8823 26970
rect 9345 26966 9348 26992
rect 9374 26966 9377 26992
rect 10734 26990 10748 27006
rect 11599 27000 11602 27006
rect 11628 27000 11631 27026
rect 11838 27024 11852 27040
rect 13255 27034 13258 27060
rect 13284 27054 13287 27060
rect 13494 27058 13508 27074
rect 16337 27068 16340 27094
rect 16366 27068 16369 27094
rect 16475 27068 16478 27094
rect 16504 27068 16507 27094
rect 13348 27055 13377 27058
rect 13348 27054 13354 27055
rect 13284 27040 13354 27054
rect 13284 27034 13287 27040
rect 13348 27038 13354 27040
rect 13371 27038 13377 27055
rect 13348 27035 13377 27038
rect 13394 27055 13423 27058
rect 13394 27038 13400 27055
rect 13417 27038 13423 27055
rect 13394 27035 13423 27038
rect 13486 27055 13515 27058
rect 13486 27038 13492 27055
rect 13509 27054 13515 27055
rect 13715 27054 13718 27060
rect 13509 27040 13718 27054
rect 13509 27038 13515 27040
rect 13486 27035 13515 27038
rect 11830 27021 11859 27024
rect 11830 27004 11836 27021
rect 11853 27004 11859 27021
rect 13402 27020 13416 27035
rect 13715 27034 13718 27040
rect 13744 27034 13747 27060
rect 14589 27034 14592 27060
rect 14618 27034 14621 27060
rect 15095 27034 15098 27060
rect 15124 27054 15127 27060
rect 16522 27055 16551 27058
rect 16522 27054 16528 27055
rect 15124 27040 16528 27054
rect 15124 27034 15127 27040
rect 16522 27038 16528 27040
rect 16545 27054 16551 27055
rect 17303 27054 17306 27060
rect 16545 27040 17306 27054
rect 16545 27038 16551 27040
rect 16522 27035 16551 27038
rect 17303 27034 17306 27040
rect 17332 27034 17335 27060
rect 18223 27034 18226 27060
rect 18252 27034 18255 27060
rect 18269 27034 18272 27060
rect 18298 27034 18301 27060
rect 18361 27034 18364 27060
rect 18390 27034 18393 27060
rect 20155 27034 20158 27060
rect 20184 27054 20187 27060
rect 20293 27054 20296 27060
rect 20184 27040 20296 27054
rect 20184 27034 20187 27040
rect 20293 27034 20296 27040
rect 20322 27034 20325 27060
rect 20431 27034 20434 27060
rect 20460 27034 20463 27060
rect 21121 27034 21124 27060
rect 21150 27054 21153 27060
rect 21306 27055 21335 27058
rect 21306 27054 21312 27055
rect 21150 27040 21312 27054
rect 21150 27034 21153 27040
rect 21306 27038 21312 27040
rect 21329 27038 21335 27055
rect 21306 27035 21335 27038
rect 13577 27020 13580 27026
rect 13402 27006 13580 27020
rect 11830 27001 11859 27004
rect 13577 27000 13580 27006
rect 13606 27000 13609 27026
rect 10726 26987 10755 26990
rect 10726 26970 10732 26987
rect 10749 26970 10755 26987
rect 10726 26967 10755 26970
rect 10817 26966 10820 26992
rect 10846 26966 10849 26992
rect 11875 26966 11878 26992
rect 11904 26986 11907 26992
rect 12198 26987 12227 26990
rect 12198 26986 12204 26987
rect 11904 26972 12204 26986
rect 11904 26966 11907 26972
rect 12198 26970 12204 26972
rect 12221 26970 12227 26987
rect 12198 26967 12227 26970
rect 16568 26987 16597 26990
rect 16568 26970 16574 26987
rect 16591 26986 16597 26987
rect 16613 26986 16616 26992
rect 16591 26972 16616 26986
rect 16591 26970 16597 26972
rect 16568 26967 16597 26970
rect 16613 26966 16616 26972
rect 16642 26966 16645 26992
rect 3036 26904 29992 26952
rect 17948 26885 17977 26888
rect 17948 26868 17954 26885
rect 17971 26884 17977 26885
rect 18269 26884 18272 26890
rect 17971 26870 18272 26884
rect 17971 26868 17977 26870
rect 17948 26865 17977 26868
rect 18269 26864 18272 26870
rect 18298 26864 18301 26890
rect 6907 26850 6910 26856
rect 6778 26836 6910 26850
rect 6778 26820 6792 26836
rect 6907 26830 6910 26836
rect 6936 26850 6939 26856
rect 7505 26850 7508 26856
rect 6936 26836 7508 26850
rect 6936 26830 6939 26836
rect 7505 26830 7508 26836
rect 7534 26830 7537 26856
rect 15049 26830 15052 26856
rect 15078 26830 15081 26856
rect 6770 26817 6799 26820
rect 6770 26800 6776 26817
rect 6793 26800 6799 26817
rect 6770 26797 6799 26800
rect 6999 26796 7002 26822
rect 7028 26816 7031 26822
rect 7598 26817 7627 26820
rect 7598 26816 7604 26817
rect 7028 26802 7604 26816
rect 7028 26796 7031 26802
rect 7598 26800 7604 26802
rect 7621 26800 7627 26817
rect 7598 26797 7627 26800
rect 7644 26817 7673 26820
rect 7644 26800 7650 26817
rect 7667 26816 7673 26817
rect 7689 26816 7692 26822
rect 7667 26802 7692 26816
rect 7667 26800 7673 26802
rect 7644 26797 7673 26800
rect 7689 26796 7692 26802
rect 7718 26816 7721 26822
rect 8195 26816 8198 26822
rect 7718 26802 8198 26816
rect 7718 26796 7721 26802
rect 8195 26796 8198 26802
rect 8224 26796 8227 26822
rect 8655 26796 8658 26822
rect 8684 26796 8687 26822
rect 13623 26796 13626 26822
rect 13652 26816 13655 26822
rect 14589 26816 14592 26822
rect 13652 26802 14592 26816
rect 13652 26796 13655 26802
rect 14589 26796 14592 26802
rect 14618 26816 14621 26822
rect 16476 26817 16505 26820
rect 16476 26816 16482 26817
rect 14618 26802 16482 26816
rect 14618 26796 14621 26802
rect 16476 26800 16482 26802
rect 16499 26800 16505 26817
rect 16476 26797 16505 26800
rect 17994 26817 18023 26820
rect 17994 26800 18000 26817
rect 18017 26816 18023 26817
rect 18453 26816 18456 26822
rect 18017 26802 18456 26816
rect 18017 26800 18023 26802
rect 17994 26797 18023 26800
rect 18453 26796 18456 26802
rect 18482 26796 18485 26822
rect 6631 26762 6634 26788
rect 6660 26762 6663 26788
rect 6861 26762 6864 26788
rect 6890 26782 6893 26788
rect 6954 26783 6983 26786
rect 6954 26782 6960 26783
rect 6890 26768 6960 26782
rect 6890 26762 6893 26768
rect 6954 26766 6960 26768
rect 6977 26766 6983 26783
rect 6954 26763 6983 26766
rect 7506 26783 7535 26786
rect 7506 26766 7512 26783
rect 7529 26766 7535 26783
rect 7506 26763 7535 26766
rect 6999 26728 7002 26754
rect 7028 26748 7031 26754
rect 7414 26749 7443 26752
rect 7414 26748 7420 26749
rect 7028 26734 7420 26748
rect 7028 26728 7031 26734
rect 7414 26732 7420 26734
rect 7437 26732 7443 26749
rect 7414 26729 7443 26732
rect 7514 26748 7528 26763
rect 7551 26762 7554 26788
rect 7580 26762 7583 26788
rect 8609 26782 8612 26788
rect 7698 26768 8612 26782
rect 7698 26748 7712 26768
rect 8609 26762 8612 26768
rect 8638 26762 8641 26788
rect 10219 26762 10222 26788
rect 10248 26782 10251 26788
rect 10266 26783 10295 26786
rect 10266 26782 10272 26783
rect 10248 26768 10272 26782
rect 10248 26762 10251 26768
rect 10266 26766 10272 26768
rect 10289 26766 10295 26783
rect 10266 26763 10295 26766
rect 10400 26783 10429 26786
rect 10400 26766 10406 26783
rect 10423 26782 10429 26783
rect 10817 26782 10820 26788
rect 10423 26768 10820 26782
rect 10423 26766 10429 26768
rect 10400 26763 10429 26766
rect 7514 26734 7712 26748
rect 8518 26749 8547 26752
rect 7275 26694 7278 26720
rect 7304 26714 7307 26720
rect 7514 26714 7528 26734
rect 8518 26732 8524 26749
rect 8541 26748 8547 26749
rect 8931 26748 8934 26754
rect 8541 26734 8934 26748
rect 8541 26732 8547 26734
rect 8518 26729 8547 26732
rect 8931 26728 8934 26734
rect 8960 26728 8963 26754
rect 10274 26748 10288 26763
rect 10817 26762 10820 26768
rect 10846 26762 10849 26788
rect 11278 26783 11307 26786
rect 11278 26766 11284 26783
rect 11301 26766 11307 26783
rect 11278 26763 11307 26766
rect 11412 26783 11441 26786
rect 11412 26766 11418 26783
rect 11435 26782 11441 26783
rect 11875 26782 11878 26788
rect 11435 26768 11878 26782
rect 11435 26766 11441 26768
rect 11412 26763 11441 26766
rect 11047 26748 11050 26754
rect 10274 26734 11050 26748
rect 11047 26728 11050 26734
rect 11076 26748 11079 26754
rect 11286 26748 11300 26763
rect 11875 26762 11878 26768
rect 11904 26762 11907 26788
rect 12197 26762 12200 26788
rect 12226 26762 12229 26788
rect 12289 26762 12292 26788
rect 12318 26762 12321 26788
rect 14636 26783 14665 26786
rect 14636 26766 14642 26783
rect 14659 26782 14665 26783
rect 14866 26783 14895 26786
rect 14866 26782 14872 26783
rect 14659 26768 14872 26782
rect 14659 26766 14665 26768
rect 14636 26763 14665 26766
rect 14866 26766 14872 26768
rect 14889 26766 14895 26783
rect 14866 26763 14895 26766
rect 14943 26783 14972 26786
rect 14943 26766 14949 26783
rect 14966 26782 14972 26783
rect 15141 26782 15144 26788
rect 14966 26768 15144 26782
rect 14966 26766 14972 26768
rect 14943 26763 14972 26766
rect 11737 26748 11740 26754
rect 11076 26734 11740 26748
rect 11076 26728 11079 26734
rect 11737 26728 11740 26734
rect 11766 26748 11769 26754
rect 13117 26748 13120 26754
rect 11766 26734 13120 26748
rect 11766 26728 11769 26734
rect 13117 26728 13120 26734
rect 13146 26748 13149 26754
rect 13623 26748 13626 26754
rect 13146 26734 13626 26748
rect 13146 26728 13149 26734
rect 13623 26728 13626 26734
rect 13652 26728 13655 26754
rect 14874 26748 14888 26763
rect 15141 26762 15144 26768
rect 15170 26762 15173 26788
rect 16613 26786 16616 26788
rect 16610 26782 16616 26786
rect 16593 26768 16616 26782
rect 16610 26763 16616 26768
rect 16613 26762 16616 26763
rect 16642 26762 16645 26788
rect 17809 26762 17812 26788
rect 17838 26762 17841 26788
rect 19097 26762 19100 26788
rect 19126 26782 19129 26788
rect 19144 26783 19173 26786
rect 19144 26782 19150 26783
rect 19126 26768 19150 26782
rect 19126 26762 19129 26768
rect 19144 26766 19150 26768
rect 19167 26766 19173 26783
rect 19144 26763 19173 26766
rect 17671 26748 17674 26754
rect 14874 26734 17674 26748
rect 17671 26728 17674 26734
rect 17700 26728 17703 26754
rect 18637 26728 18640 26754
rect 18666 26748 18669 26754
rect 19373 26752 19376 26754
rect 19304 26749 19333 26752
rect 19304 26748 19310 26749
rect 18666 26734 19310 26748
rect 18666 26728 18669 26734
rect 19304 26732 19310 26734
rect 19327 26732 19333 26749
rect 19304 26729 19333 26732
rect 19355 26749 19376 26752
rect 19355 26732 19361 26749
rect 19355 26729 19376 26732
rect 19373 26728 19376 26729
rect 19402 26728 19405 26754
rect 7304 26700 7528 26714
rect 8334 26715 8363 26718
rect 7304 26694 7307 26700
rect 8334 26698 8340 26715
rect 8357 26714 8363 26715
rect 8471 26714 8474 26720
rect 8357 26700 8474 26714
rect 8357 26698 8363 26700
rect 8334 26695 8363 26698
rect 8471 26694 8474 26700
rect 8500 26694 8503 26720
rect 8563 26694 8566 26720
rect 8592 26694 8595 26720
rect 10541 26694 10544 26720
rect 10570 26714 10573 26720
rect 10956 26715 10985 26718
rect 10956 26714 10962 26715
rect 10570 26700 10962 26714
rect 10570 26694 10573 26700
rect 10956 26698 10962 26700
rect 10979 26698 10985 26715
rect 10956 26695 10985 26698
rect 11967 26694 11970 26720
rect 11996 26694 11999 26720
rect 12243 26694 12246 26720
rect 12272 26694 12275 26720
rect 17165 26694 17168 26720
rect 17194 26694 17197 26720
rect 17763 26694 17766 26720
rect 17792 26714 17795 26720
rect 17856 26715 17885 26718
rect 17856 26714 17862 26715
rect 17792 26700 17862 26714
rect 17792 26694 17795 26700
rect 17856 26698 17862 26700
rect 17879 26698 17885 26715
rect 17856 26695 17885 26698
rect 17901 26694 17904 26720
rect 17930 26694 17933 26720
rect 20179 26715 20208 26718
rect 20179 26698 20185 26715
rect 20202 26714 20208 26715
rect 20615 26714 20618 26720
rect 20202 26700 20618 26714
rect 20202 26698 20208 26700
rect 20179 26695 20208 26698
rect 20615 26694 20618 26700
rect 20644 26694 20647 26720
rect 3036 26632 29992 26680
rect 6217 26592 6220 26618
rect 6246 26612 6249 26618
rect 6264 26613 6293 26616
rect 6264 26612 6270 26613
rect 6246 26598 6270 26612
rect 6246 26592 6249 26598
rect 6264 26596 6270 26598
rect 6287 26596 6293 26613
rect 6264 26593 6293 26596
rect 6631 26592 6634 26618
rect 6660 26612 6663 26618
rect 6954 26613 6983 26616
rect 6954 26612 6960 26613
rect 6660 26598 6960 26612
rect 6660 26592 6663 26598
rect 6954 26596 6960 26598
rect 6977 26596 6983 26613
rect 6954 26593 6983 26596
rect 7183 26592 7186 26618
rect 7212 26612 7215 26618
rect 7551 26612 7554 26618
rect 7212 26598 7554 26612
rect 7212 26592 7215 26598
rect 7551 26592 7554 26598
rect 7580 26592 7583 26618
rect 10725 26592 10728 26618
rect 10754 26592 10757 26618
rect 17395 26612 17398 26618
rect 15794 26598 17398 26612
rect 6217 26524 6220 26550
rect 6246 26524 6249 26550
rect 6264 26511 6293 26514
rect 6264 26494 6270 26511
rect 6287 26494 6293 26511
rect 6264 26491 6293 26494
rect 6356 26511 6385 26514
rect 6356 26494 6362 26511
rect 6379 26510 6385 26511
rect 6640 26510 6654 26592
rect 7689 26578 7692 26584
rect 7146 26564 7692 26578
rect 6953 26524 6956 26550
rect 6982 26524 6985 26550
rect 7046 26545 7075 26548
rect 7046 26528 7052 26545
rect 7069 26544 7075 26545
rect 7146 26544 7160 26564
rect 7689 26558 7692 26564
rect 7718 26558 7721 26584
rect 11872 26579 11901 26582
rect 11872 26562 11878 26579
rect 11895 26578 11901 26579
rect 12243 26578 12246 26584
rect 11895 26564 12246 26578
rect 11895 26562 11901 26564
rect 11872 26559 11901 26562
rect 12243 26558 12246 26564
rect 12272 26558 12275 26584
rect 15794 26582 15808 26598
rect 17395 26592 17398 26598
rect 17424 26612 17427 26618
rect 17809 26612 17812 26618
rect 17424 26598 17812 26612
rect 17424 26592 17427 26598
rect 17809 26592 17812 26598
rect 17838 26592 17841 26618
rect 20386 26613 20415 26616
rect 20386 26596 20392 26613
rect 20409 26612 20415 26613
rect 20431 26612 20434 26618
rect 20409 26598 20434 26612
rect 20409 26596 20415 26598
rect 20386 26593 20415 26596
rect 20431 26592 20434 26598
rect 20460 26592 20463 26618
rect 20615 26592 20618 26618
rect 20644 26592 20647 26618
rect 15786 26579 15815 26582
rect 15786 26562 15792 26579
rect 15809 26562 15815 26579
rect 15786 26559 15815 26562
rect 15831 26558 15834 26584
rect 15860 26578 15863 26584
rect 15878 26579 15907 26582
rect 15878 26578 15884 26579
rect 15860 26564 15884 26578
rect 15860 26558 15863 26564
rect 15878 26562 15884 26564
rect 15901 26562 15907 26579
rect 17211 26578 17214 26584
rect 15878 26559 15907 26562
rect 16254 26564 17214 26578
rect 7069 26530 7160 26544
rect 7069 26528 7075 26530
rect 7046 26525 7075 26528
rect 7183 26524 7186 26550
rect 7212 26524 7215 26550
rect 7275 26524 7278 26550
rect 7304 26524 7307 26550
rect 9253 26524 9256 26550
rect 9282 26524 9285 26550
rect 10541 26524 10544 26550
rect 10570 26524 10573 26550
rect 11737 26524 11740 26550
rect 11766 26524 11769 26550
rect 13485 26524 13488 26550
rect 13514 26524 13517 26550
rect 13531 26524 13534 26550
rect 13560 26524 13563 26550
rect 13670 26545 13699 26548
rect 13670 26528 13676 26545
rect 13693 26544 13699 26545
rect 13761 26544 13764 26550
rect 13693 26530 13764 26544
rect 13693 26528 13699 26530
rect 13670 26525 13699 26528
rect 13761 26524 13764 26530
rect 13790 26524 13793 26550
rect 15188 26545 15217 26548
rect 15188 26528 15194 26545
rect 15211 26528 15217 26545
rect 15188 26525 15217 26528
rect 6379 26496 6654 26510
rect 6379 26494 6385 26496
rect 6356 26491 6385 26494
rect 6272 26476 6286 26491
rect 6861 26490 6864 26516
rect 6890 26510 6893 26516
rect 9299 26510 9302 26516
rect 6890 26496 9302 26510
rect 6890 26490 6893 26496
rect 9299 26490 9302 26496
rect 9328 26490 9331 26516
rect 9345 26490 9348 26516
rect 9374 26490 9377 26516
rect 10495 26490 10498 26516
rect 10524 26490 10527 26516
rect 13577 26490 13580 26516
rect 13606 26490 13609 26516
rect 14957 26490 14960 26516
rect 14986 26510 14989 26516
rect 15142 26511 15171 26514
rect 15142 26510 15148 26511
rect 14986 26496 15148 26510
rect 14986 26490 14989 26496
rect 15142 26494 15148 26496
rect 15165 26494 15171 26511
rect 15142 26491 15171 26494
rect 6870 26476 6884 26490
rect 6272 26462 6884 26476
rect 15196 26476 15210 26525
rect 15923 26524 15926 26550
rect 15952 26524 15955 26550
rect 16254 26548 16268 26564
rect 17211 26558 17214 26564
rect 17240 26578 17243 26584
rect 20570 26579 20599 26582
rect 17240 26564 18338 26578
rect 17240 26558 17243 26564
rect 16246 26545 16275 26548
rect 16246 26528 16252 26545
rect 16269 26528 16275 26545
rect 16246 26525 16275 26528
rect 17165 26524 17168 26550
rect 17194 26544 17197 26550
rect 17810 26545 17839 26548
rect 17810 26544 17816 26545
rect 17194 26530 17816 26544
rect 17194 26524 17197 26530
rect 17810 26528 17816 26530
rect 17833 26528 17839 26545
rect 17810 26525 17839 26528
rect 18039 26524 18042 26550
rect 18068 26544 18071 26550
rect 18324 26548 18338 26564
rect 20570 26562 20576 26579
rect 20593 26578 20599 26579
rect 21121 26578 21124 26584
rect 20593 26564 21124 26578
rect 20593 26562 20599 26564
rect 20570 26559 20599 26562
rect 21121 26558 21124 26564
rect 21150 26558 21153 26584
rect 21283 26579 21312 26582
rect 21283 26578 21289 26579
rect 21176 26564 21289 26578
rect 18224 26545 18253 26548
rect 18224 26544 18230 26545
rect 18068 26530 18230 26544
rect 18068 26524 18071 26530
rect 18224 26528 18230 26530
rect 18247 26528 18253 26545
rect 18224 26525 18253 26528
rect 18316 26545 18345 26548
rect 18316 26528 18322 26545
rect 18339 26544 18345 26545
rect 18499 26544 18502 26550
rect 18339 26530 18502 26544
rect 18339 26528 18345 26530
rect 18316 26525 18345 26528
rect 18499 26524 18502 26530
rect 18528 26524 18531 26550
rect 20247 26524 20250 26550
rect 20276 26544 20279 26550
rect 21176 26544 21190 26564
rect 21283 26562 21289 26564
rect 21306 26562 21312 26579
rect 21283 26559 21312 26562
rect 20276 26530 21190 26544
rect 21237 26545 21266 26548
rect 20276 26524 20279 26530
rect 21237 26528 21243 26545
rect 21260 26544 21266 26545
rect 21489 26544 21492 26550
rect 21260 26530 21492 26544
rect 21260 26528 21266 26530
rect 21237 26525 21266 26528
rect 21489 26524 21492 26530
rect 21518 26524 21521 26550
rect 15372 26511 15401 26514
rect 15372 26494 15378 26511
rect 15395 26510 15401 26511
rect 16200 26511 16229 26514
rect 16200 26510 16206 26511
rect 15395 26496 16206 26510
rect 15395 26494 15401 26496
rect 15372 26491 15401 26494
rect 16200 26494 16206 26496
rect 16223 26510 16229 26511
rect 16337 26510 16340 26516
rect 16223 26496 16340 26510
rect 16223 26494 16229 26496
rect 16200 26491 16229 26494
rect 16337 26490 16340 26496
rect 16366 26490 16369 26516
rect 17174 26476 17188 26524
rect 17717 26490 17720 26516
rect 17746 26510 17749 26516
rect 17764 26511 17793 26514
rect 17764 26510 17770 26511
rect 17746 26496 17770 26510
rect 17746 26490 17749 26496
rect 17764 26494 17770 26496
rect 17787 26494 17793 26511
rect 17764 26491 17793 26494
rect 17901 26490 17904 26516
rect 17930 26510 17933 26516
rect 17994 26511 18023 26514
rect 17994 26510 18000 26511
rect 17930 26496 18000 26510
rect 17930 26490 17933 26496
rect 17994 26494 18000 26496
rect 18017 26494 18023 26511
rect 17994 26491 18023 26494
rect 20661 26490 20664 26516
rect 20690 26490 20693 26516
rect 21076 26511 21105 26514
rect 21076 26494 21082 26511
rect 21099 26494 21105 26511
rect 21076 26491 21105 26494
rect 18224 26477 18253 26480
rect 18224 26476 18230 26477
rect 15196 26462 17188 26476
rect 17933 26462 18230 26476
rect 5849 26422 5852 26448
rect 5878 26442 5881 26448
rect 6034 26443 6063 26446
rect 6034 26442 6040 26443
rect 5878 26428 6040 26442
rect 5878 26422 5881 26428
rect 6034 26426 6040 26428
rect 6057 26426 6063 26443
rect 6034 26423 6063 26426
rect 9069 26422 9072 26448
rect 9098 26422 9101 26448
rect 12428 26443 12457 26446
rect 12428 26426 12434 26443
rect 12451 26442 12457 26443
rect 12473 26442 12476 26448
rect 12451 26428 12476 26442
rect 12451 26426 12457 26428
rect 12428 26423 12457 26426
rect 12473 26422 12476 26428
rect 12502 26422 12505 26448
rect 13669 26422 13672 26448
rect 13698 26422 13701 26448
rect 15924 26443 15953 26446
rect 15924 26426 15930 26443
rect 15947 26442 15953 26443
rect 16199 26442 16202 26448
rect 15947 26428 16202 26442
rect 15947 26426 15953 26428
rect 15924 26423 15953 26426
rect 16199 26422 16202 26428
rect 16228 26422 16231 26448
rect 16337 26422 16340 26448
rect 16366 26442 16369 26448
rect 16384 26443 16413 26446
rect 16384 26442 16390 26443
rect 16366 26428 16390 26442
rect 16366 26422 16369 26428
rect 16384 26426 16390 26428
rect 16407 26426 16413 26443
rect 16384 26423 16413 26426
rect 17855 26422 17858 26448
rect 17884 26442 17887 26448
rect 17933 26442 17947 26462
rect 18224 26460 18230 26462
rect 18247 26460 18253 26477
rect 18224 26457 18253 26460
rect 19097 26456 19100 26482
rect 19126 26476 19129 26482
rect 20293 26476 20296 26482
rect 19126 26462 20296 26476
rect 19126 26456 19129 26462
rect 20293 26456 20296 26462
rect 20322 26476 20325 26482
rect 21084 26476 21098 26491
rect 20322 26462 21098 26476
rect 20322 26456 20325 26462
rect 22133 26446 22136 26448
rect 17884 26428 17947 26442
rect 22111 26443 22136 26446
rect 17884 26422 17887 26428
rect 22111 26426 22117 26443
rect 22134 26426 22136 26443
rect 22111 26423 22136 26426
rect 22133 26422 22136 26423
rect 22162 26422 22165 26448
rect 3036 26360 29992 26408
rect 6217 26320 6220 26346
rect 6246 26340 6249 26346
rect 6563 26341 6592 26344
rect 6563 26340 6569 26341
rect 6246 26326 6569 26340
rect 6246 26320 6249 26326
rect 6563 26324 6569 26326
rect 6586 26324 6592 26341
rect 6563 26321 6592 26324
rect 7505 26320 7508 26346
rect 7534 26340 7537 26346
rect 8563 26340 8566 26346
rect 7534 26326 8566 26340
rect 7534 26320 7537 26326
rect 8020 26276 8034 26326
rect 8563 26320 8566 26326
rect 8592 26320 8595 26346
rect 12106 26341 12135 26344
rect 12106 26324 12112 26341
rect 12129 26340 12135 26341
rect 12197 26340 12200 26346
rect 12129 26326 12200 26340
rect 12129 26324 12135 26326
rect 12106 26321 12135 26324
rect 12197 26320 12200 26326
rect 12226 26320 12229 26346
rect 13103 26326 14244 26340
rect 10817 26286 10820 26312
rect 10846 26306 10849 26312
rect 13103 26306 13117 26326
rect 10846 26292 13117 26306
rect 14230 26306 14244 26326
rect 16337 26320 16340 26346
rect 16366 26320 16369 26346
rect 17855 26320 17858 26346
rect 17884 26320 17887 26346
rect 17257 26306 17260 26312
rect 14230 26292 17260 26306
rect 10846 26286 10849 26292
rect 17257 26286 17260 26292
rect 17286 26286 17289 26312
rect 17993 26286 17996 26312
rect 18022 26306 18025 26312
rect 18022 26292 19120 26306
rect 18022 26286 18025 26292
rect 8012 26273 8041 26276
rect 8012 26256 8018 26273
rect 8035 26256 8041 26273
rect 8012 26253 8041 26256
rect 8104 26273 8133 26276
rect 8104 26256 8110 26273
rect 8127 26272 8133 26273
rect 8333 26272 8336 26278
rect 8127 26258 8336 26272
rect 8127 26256 8133 26258
rect 8104 26253 8133 26256
rect 8333 26252 8336 26258
rect 8362 26252 8365 26278
rect 9299 26252 9302 26278
rect 9328 26272 9331 26278
rect 13302 26273 13331 26276
rect 9328 26258 13094 26272
rect 9328 26252 9331 26258
rect 5527 26218 5530 26244
rect 5556 26218 5559 26244
rect 5689 26239 5718 26242
rect 5689 26222 5695 26239
rect 5712 26238 5718 26239
rect 5849 26238 5852 26244
rect 5712 26224 5852 26238
rect 5712 26222 5718 26224
rect 5689 26219 5718 26222
rect 5849 26218 5852 26224
rect 5878 26218 5881 26244
rect 8425 26218 8428 26244
rect 8454 26218 8457 26244
rect 8471 26218 8474 26244
rect 8500 26238 8503 26244
rect 8581 26239 8610 26242
rect 8581 26238 8587 26239
rect 8500 26224 8587 26238
rect 8500 26218 8503 26224
rect 8581 26222 8587 26224
rect 8604 26222 8610 26239
rect 8581 26219 8610 26222
rect 11599 26218 11602 26244
rect 11628 26218 11631 26244
rect 11700 26242 11714 26258
rect 11692 26239 11721 26242
rect 11692 26222 11698 26239
rect 11715 26222 11721 26239
rect 11692 26219 11721 26222
rect 12106 26239 12135 26242
rect 12106 26222 12112 26239
rect 12129 26222 12135 26239
rect 12106 26219 12135 26222
rect 12198 26239 12227 26242
rect 12198 26222 12204 26239
rect 12221 26238 12227 26239
rect 12473 26238 12476 26244
rect 12221 26224 12476 26238
rect 12221 26222 12227 26224
rect 12198 26219 12227 26222
rect 5573 26184 5576 26210
rect 5602 26204 5605 26210
rect 5735 26205 5764 26208
rect 5735 26204 5741 26205
rect 5602 26190 5741 26204
rect 5602 26184 5605 26190
rect 5735 26188 5741 26190
rect 5758 26188 5764 26205
rect 5735 26185 5764 26188
rect 6769 26184 6772 26210
rect 6798 26204 6801 26210
rect 7505 26204 7508 26210
rect 6798 26190 7508 26204
rect 6798 26184 6801 26190
rect 7505 26184 7508 26190
rect 7534 26204 7537 26210
rect 7966 26205 7995 26208
rect 7534 26190 7942 26204
rect 7534 26184 7537 26190
rect 6563 26171 6592 26174
rect 6563 26154 6569 26171
rect 6586 26170 6592 26171
rect 7229 26170 7232 26176
rect 6586 26156 7232 26170
rect 6586 26154 6592 26156
rect 6563 26151 6592 26154
rect 7229 26150 7232 26156
rect 7258 26150 7261 26176
rect 7551 26150 7554 26176
rect 7580 26170 7583 26176
rect 7782 26171 7811 26174
rect 7782 26170 7788 26171
rect 7580 26156 7788 26170
rect 7580 26150 7583 26156
rect 7782 26154 7788 26156
rect 7805 26154 7811 26171
rect 7928 26170 7942 26190
rect 7966 26188 7972 26205
rect 7989 26204 7995 26205
rect 8241 26204 8244 26210
rect 7989 26190 8244 26204
rect 7989 26188 7995 26190
rect 7966 26185 7995 26188
rect 8241 26184 8244 26190
rect 8270 26184 8273 26210
rect 8625 26205 8654 26208
rect 8625 26204 8631 26205
rect 8296 26190 8631 26204
rect 8296 26170 8310 26190
rect 8625 26188 8631 26190
rect 8648 26204 8654 26205
rect 8701 26204 8704 26210
rect 8648 26190 8704 26204
rect 8648 26188 8654 26190
rect 8625 26185 8654 26188
rect 8701 26184 8704 26190
rect 8730 26184 8733 26210
rect 11646 26205 11675 26208
rect 11646 26188 11652 26205
rect 11669 26204 11675 26205
rect 12114 26204 12128 26219
rect 12473 26218 12476 26224
rect 12502 26218 12505 26244
rect 12934 26239 12963 26242
rect 12934 26222 12940 26239
rect 12957 26238 12963 26239
rect 13025 26238 13028 26244
rect 12957 26224 13028 26238
rect 12957 26222 12963 26224
rect 12934 26219 12963 26222
rect 13025 26218 13028 26224
rect 13054 26218 13057 26244
rect 13080 26238 13094 26258
rect 13302 26256 13308 26273
rect 13325 26272 13331 26273
rect 13531 26272 13534 26278
rect 13325 26258 13534 26272
rect 13325 26256 13331 26258
rect 13302 26253 13331 26256
rect 13531 26252 13534 26258
rect 13560 26252 13563 26278
rect 13623 26252 13626 26278
rect 13652 26252 13655 26278
rect 14451 26252 14454 26278
rect 14480 26272 14483 26278
rect 14480 26258 14842 26272
rect 14480 26252 14483 26258
rect 13080 26224 13232 26238
rect 11669 26190 12128 26204
rect 13218 26204 13232 26224
rect 13255 26218 13258 26244
rect 13284 26218 13287 26244
rect 13310 26224 13646 26238
rect 13310 26204 13324 26224
rect 13218 26190 13324 26204
rect 13632 26204 13646 26224
rect 13669 26218 13672 26244
rect 13698 26238 13701 26244
rect 13752 26239 13781 26242
rect 13752 26238 13758 26239
rect 13698 26224 13758 26238
rect 13698 26218 13701 26224
rect 13752 26222 13758 26224
rect 13775 26222 13781 26239
rect 14129 26238 14132 26244
rect 13752 26219 13781 26222
rect 13816 26224 14132 26238
rect 13816 26204 13830 26224
rect 14129 26218 14132 26224
rect 14158 26218 14161 26244
rect 14774 26239 14803 26242
rect 14774 26238 14780 26239
rect 14184 26224 14780 26238
rect 14184 26204 14198 26224
rect 14774 26222 14780 26224
rect 14797 26222 14803 26239
rect 14828 26238 14842 26258
rect 14957 26252 14960 26278
rect 14986 26252 14989 26278
rect 18867 26272 18870 26278
rect 16346 26258 18870 26272
rect 15050 26239 15079 26242
rect 15050 26238 15056 26239
rect 14828 26224 15056 26238
rect 14774 26219 14803 26222
rect 15050 26222 15056 26224
rect 15073 26222 15079 26239
rect 15050 26219 15079 26222
rect 16291 26218 16294 26244
rect 16320 26218 16323 26244
rect 16346 26242 16360 26258
rect 18867 26252 18870 26258
rect 18896 26252 18899 26278
rect 19106 26272 19120 26292
rect 19106 26258 19166 26272
rect 16338 26239 16367 26242
rect 16338 26222 16344 26239
rect 16361 26222 16367 26239
rect 16338 26219 16367 26222
rect 17303 26218 17306 26244
rect 17332 26238 17335 26244
rect 17902 26239 17931 26242
rect 17902 26238 17908 26239
rect 17332 26224 17908 26238
rect 17332 26218 17335 26224
rect 17902 26222 17908 26224
rect 17925 26222 17931 26239
rect 17902 26219 17931 26222
rect 19097 26218 19100 26244
rect 19126 26218 19129 26244
rect 19152 26238 19166 26258
rect 19373 26238 19376 26244
rect 19152 26224 19376 26238
rect 13632 26190 13830 26204
rect 14138 26190 14198 26204
rect 11669 26188 11675 26190
rect 11646 26185 11675 26188
rect 7928 26156 8310 26170
rect 7782 26151 7811 26154
rect 8931 26150 8934 26176
rect 8960 26170 8963 26176
rect 9461 26171 9490 26174
rect 9461 26170 9467 26171
rect 8960 26156 9467 26170
rect 8960 26150 8963 26156
rect 9461 26154 9467 26156
rect 9484 26154 9490 26171
rect 9461 26151 9490 26154
rect 13255 26150 13258 26176
rect 13284 26170 13287 26176
rect 14138 26170 14152 26190
rect 16199 26184 16202 26210
rect 16228 26184 16231 26210
rect 17487 26184 17490 26210
rect 17516 26204 17519 26210
rect 17717 26204 17720 26210
rect 17516 26190 17720 26204
rect 17516 26184 17519 26190
rect 17717 26184 17720 26190
rect 17746 26184 17749 26210
rect 17947 26184 17950 26210
rect 17976 26184 17979 26210
rect 18637 26184 18640 26210
rect 18666 26204 18669 26210
rect 19313 26208 19327 26224
rect 19373 26218 19376 26224
rect 19402 26218 19405 26244
rect 19258 26205 19287 26208
rect 19258 26204 19264 26205
rect 18666 26190 19264 26204
rect 18666 26184 18669 26190
rect 19258 26188 19264 26190
rect 19281 26188 19287 26205
rect 19258 26185 19287 26188
rect 19305 26205 19334 26208
rect 19305 26188 19311 26205
rect 19328 26188 19334 26205
rect 19305 26185 19334 26188
rect 20133 26205 20162 26208
rect 20133 26188 20139 26205
rect 20156 26204 20162 26205
rect 20523 26204 20526 26210
rect 20156 26190 20526 26204
rect 20156 26188 20162 26190
rect 20133 26185 20162 26188
rect 20523 26184 20526 26190
rect 20552 26184 20555 26210
rect 13284 26156 14152 26170
rect 14314 26171 14343 26174
rect 13284 26150 13287 26156
rect 14314 26154 14320 26171
rect 14337 26170 14343 26171
rect 14451 26170 14454 26176
rect 14337 26156 14454 26170
rect 14337 26154 14343 26156
rect 14314 26151 14343 26154
rect 14451 26150 14454 26156
rect 14480 26150 14483 26176
rect 16429 26150 16432 26176
rect 16458 26150 16461 26176
rect 17671 26150 17674 26176
rect 17700 26170 17703 26176
rect 17764 26171 17793 26174
rect 17764 26170 17770 26171
rect 17700 26156 17770 26170
rect 17700 26150 17703 26156
rect 17764 26154 17770 26156
rect 17787 26170 17793 26171
rect 17993 26170 17996 26176
rect 17787 26156 17996 26170
rect 17787 26154 17793 26156
rect 17764 26151 17793 26154
rect 17993 26150 17996 26156
rect 18022 26150 18025 26176
rect 3036 26088 29992 26136
rect 6907 26048 6910 26074
rect 6936 26048 6939 26074
rect 13761 26048 13764 26074
rect 13790 26048 13793 26074
rect 18499 26048 18502 26074
rect 18528 26048 18531 26074
rect 4469 26014 4472 26040
rect 4498 26034 4501 26040
rect 7505 26038 7508 26040
rect 4631 26035 4660 26038
rect 4631 26034 4637 26035
rect 4498 26020 4637 26034
rect 4498 26014 4501 26020
rect 4631 26018 4637 26020
rect 4654 26018 4660 26035
rect 4631 26015 4660 26018
rect 7487 26035 7508 26038
rect 7487 26018 7493 26035
rect 7487 26015 7508 26018
rect 7505 26014 7508 26015
rect 7534 26014 7537 26040
rect 9069 26014 9072 26040
rect 9098 26034 9101 26040
rect 17947 26038 17950 26040
rect 9230 26035 9259 26038
rect 9230 26034 9236 26035
rect 9098 26020 9236 26034
rect 9098 26014 9101 26020
rect 9230 26018 9236 26020
rect 9253 26018 9259 26035
rect 9230 26015 9259 26018
rect 17944 26015 17950 26038
rect 17976 26034 17979 26040
rect 17976 26020 17994 26034
rect 17947 26014 17950 26015
rect 17976 26014 17979 26020
rect 20247 26014 20250 26040
rect 20276 26034 20279 26040
rect 20409 26035 20438 26038
rect 20409 26034 20415 26035
rect 20276 26020 20415 26034
rect 20276 26014 20279 26020
rect 20409 26018 20415 26020
rect 20432 26018 20438 26035
rect 20409 26015 20438 26018
rect 21490 26035 21519 26038
rect 21490 26018 21496 26035
rect 21513 26034 21519 26035
rect 22133 26034 22136 26040
rect 21513 26020 22136 26034
rect 21513 26018 21519 26020
rect 21490 26015 21519 26018
rect 22133 26014 22136 26020
rect 22162 26034 22165 26040
rect 23238 26035 23267 26038
rect 23238 26034 23244 26035
rect 22162 26020 23244 26034
rect 22162 26014 22165 26020
rect 23238 26018 23244 26020
rect 23261 26018 23267 26035
rect 23238 26015 23267 26018
rect 4585 26001 4614 26004
rect 4585 25984 4591 26001
rect 4608 26000 4614 26001
rect 4837 26000 4840 26006
rect 4608 25986 4840 26000
rect 4608 25984 4614 25986
rect 4585 25981 4614 25984
rect 4837 25980 4840 25986
rect 4866 26000 4869 26006
rect 6862 26001 6891 26004
rect 6862 26000 6868 26001
rect 4866 25986 6868 26000
rect 4866 25980 4869 25986
rect 6862 25984 6868 25986
rect 6885 26000 6891 26001
rect 7045 26000 7048 26006
rect 6885 25986 7048 26000
rect 6885 25984 6891 25986
rect 6862 25981 6891 25984
rect 7045 25980 7048 25986
rect 7074 25980 7077 26006
rect 7437 26001 7466 26004
rect 7437 25984 7443 26001
rect 7460 26000 7466 26001
rect 7551 26000 7554 26006
rect 7460 25986 7554 26000
rect 7460 25984 7466 25986
rect 7437 25981 7466 25984
rect 7551 25980 7554 25986
rect 7580 25980 7583 26006
rect 8701 25980 8704 26006
rect 8730 26000 8733 26006
rect 9269 26001 9298 26004
rect 9269 26000 9275 26001
rect 8730 25986 9275 26000
rect 8730 25980 8733 25986
rect 9269 25984 9275 25986
rect 9292 25984 9298 26001
rect 9269 25981 9298 25984
rect 12934 26001 12963 26004
rect 12934 25984 12940 26001
rect 12957 25984 12963 26001
rect 12934 25981 12963 25984
rect 4424 25967 4453 25970
rect 4424 25950 4430 25967
rect 4447 25950 4453 25967
rect 4424 25947 4453 25950
rect 4432 25898 4446 25947
rect 6999 25946 7002 25972
rect 7028 25946 7031 25972
rect 7276 25967 7305 25970
rect 7276 25950 7282 25967
rect 7299 25950 7305 25967
rect 7276 25947 7305 25950
rect 5527 25912 5530 25938
rect 5556 25932 5559 25938
rect 7284 25932 7298 25947
rect 8425 25946 8428 25972
rect 8454 25966 8457 25972
rect 8839 25966 8842 25972
rect 8454 25952 8842 25966
rect 8454 25946 8457 25952
rect 8839 25946 8842 25952
rect 8868 25966 8871 25972
rect 9070 25967 9099 25970
rect 9070 25966 9076 25967
rect 8868 25952 9076 25966
rect 8868 25946 8871 25952
rect 9070 25950 9076 25952
rect 9093 25950 9099 25967
rect 9070 25947 9099 25950
rect 5556 25918 7298 25932
rect 12942 25932 12956 25981
rect 13025 25980 13028 26006
rect 13054 26000 13057 26006
rect 13256 26001 13285 26004
rect 13256 26000 13262 26001
rect 13054 25986 13262 26000
rect 13054 25980 13057 25986
rect 13256 25984 13262 25986
rect 13279 25984 13285 26001
rect 13256 25981 13285 25984
rect 13394 26001 13423 26004
rect 13394 25984 13400 26001
rect 13417 26000 13423 26001
rect 13624 26001 13653 26004
rect 13624 26000 13630 26001
rect 13417 25986 13630 26000
rect 13417 25984 13423 25986
rect 13394 25981 13423 25984
rect 13624 25984 13630 25986
rect 13647 26000 13653 26001
rect 14451 26000 14454 26006
rect 13647 25986 14454 26000
rect 13647 25984 13653 25986
rect 13624 25981 13653 25984
rect 14451 25980 14454 25986
rect 14480 25980 14483 26006
rect 17810 26001 17839 26004
rect 17810 25984 17816 26001
rect 17833 26000 17839 26001
rect 20363 26001 20392 26004
rect 17833 25986 18522 26000
rect 17833 25984 17839 25986
rect 17810 25981 17839 25984
rect 18508 25972 18522 25986
rect 20363 25984 20369 26001
rect 20386 26000 20392 26001
rect 20477 26000 20480 26006
rect 20386 25986 20480 26000
rect 20386 25984 20392 25986
rect 20363 25981 20392 25984
rect 20477 25980 20480 25986
rect 20506 25980 20509 26006
rect 21351 25980 21354 26006
rect 21380 26000 21383 26006
rect 21674 26001 21703 26004
rect 21674 26000 21680 26001
rect 21380 25986 21680 26000
rect 21380 25980 21383 25986
rect 21674 25984 21680 25986
rect 21697 25984 21703 26001
rect 21674 25981 21703 25984
rect 23007 25980 23010 26006
rect 23036 26000 23039 26006
rect 23100 26001 23129 26004
rect 23100 26000 23106 26001
rect 23036 25986 23106 26000
rect 23036 25980 23039 25986
rect 23100 25984 23106 25986
rect 23123 25984 23129 26001
rect 23100 25981 23129 25984
rect 23146 26001 23175 26004
rect 23146 25984 23152 26001
rect 23169 25984 23175 26001
rect 23146 25981 23175 25984
rect 13577 25946 13580 25972
rect 13606 25966 13609 25972
rect 13670 25967 13699 25970
rect 13670 25966 13676 25967
rect 13606 25952 13676 25966
rect 13606 25946 13609 25952
rect 13670 25950 13676 25952
rect 13693 25950 13699 25967
rect 13670 25947 13699 25950
rect 13117 25932 13120 25938
rect 12942 25918 13120 25932
rect 5556 25912 5559 25918
rect 13117 25912 13120 25918
rect 13146 25932 13149 25938
rect 13255 25932 13258 25938
rect 13146 25918 13258 25932
rect 13146 25912 13149 25918
rect 13255 25912 13258 25918
rect 13284 25912 13287 25938
rect 13678 25932 13692 25947
rect 13715 25946 13718 25972
rect 13744 25966 13747 25972
rect 13762 25967 13791 25970
rect 13762 25966 13768 25967
rect 13744 25952 13768 25966
rect 13744 25946 13747 25952
rect 13762 25950 13768 25952
rect 13785 25950 13791 25967
rect 13762 25947 13791 25950
rect 18499 25946 18502 25972
rect 18528 25966 18531 25972
rect 19097 25966 19100 25972
rect 18528 25952 19100 25966
rect 18528 25946 18531 25952
rect 19097 25946 19100 25952
rect 19126 25966 19129 25972
rect 20202 25967 20231 25970
rect 20202 25966 20208 25967
rect 19126 25952 20208 25966
rect 19126 25946 19129 25952
rect 20202 25950 20208 25952
rect 20225 25950 20231 25967
rect 20202 25947 20231 25950
rect 21075 25946 21078 25972
rect 21104 25966 21107 25972
rect 21525 25967 21554 25970
rect 21525 25966 21531 25967
rect 21104 25952 21531 25966
rect 21104 25946 21107 25952
rect 21525 25950 21531 25952
rect 21548 25950 21554 25967
rect 21525 25947 21554 25950
rect 21581 25946 21584 25972
rect 21610 25966 21613 25972
rect 23154 25966 23168 25981
rect 23283 25980 23286 26006
rect 23312 25980 23315 26006
rect 23329 25980 23332 26006
rect 23358 25980 23361 26006
rect 21610 25952 23168 25966
rect 21610 25946 21613 25952
rect 23375 25946 23378 25972
rect 23404 25946 23407 25972
rect 15003 25932 15006 25938
rect 13678 25918 15006 25932
rect 15003 25912 15006 25918
rect 15032 25912 15035 25938
rect 21544 25918 21650 25932
rect 4515 25898 4518 25904
rect 4432 25884 4518 25898
rect 4515 25878 4518 25884
rect 4544 25898 4547 25904
rect 4699 25898 4702 25904
rect 4544 25884 4702 25898
rect 4544 25878 4547 25884
rect 4699 25878 4702 25884
rect 4728 25878 4731 25904
rect 5459 25899 5488 25902
rect 5459 25882 5465 25899
rect 5482 25898 5488 25899
rect 6079 25898 6082 25904
rect 5482 25884 6082 25898
rect 5482 25882 5488 25884
rect 5459 25879 5488 25882
rect 6079 25878 6082 25884
rect 6108 25878 6111 25904
rect 6631 25878 6634 25904
rect 6660 25898 6663 25904
rect 6678 25899 6707 25902
rect 6678 25898 6684 25899
rect 6660 25884 6684 25898
rect 6660 25878 6663 25884
rect 6678 25882 6684 25884
rect 6701 25882 6707 25899
rect 6678 25879 6707 25882
rect 8241 25878 8244 25904
rect 8270 25898 8273 25904
rect 8311 25899 8340 25902
rect 8311 25898 8317 25899
rect 8270 25884 8317 25898
rect 8270 25878 8273 25884
rect 8311 25882 8317 25884
rect 8334 25882 8340 25899
rect 8311 25879 8340 25882
rect 9253 25878 9256 25904
rect 9282 25898 9285 25904
rect 10127 25902 10130 25904
rect 10105 25899 10130 25902
rect 10105 25898 10111 25899
rect 9282 25884 10111 25898
rect 9282 25878 9285 25884
rect 10105 25882 10111 25884
rect 10128 25882 10130 25899
rect 10105 25879 10130 25882
rect 10127 25878 10130 25879
rect 10156 25878 10159 25904
rect 12979 25878 12982 25904
rect 13008 25898 13011 25904
rect 13072 25899 13101 25902
rect 13072 25898 13078 25899
rect 13008 25884 13078 25898
rect 13008 25878 13011 25884
rect 13072 25882 13078 25884
rect 13095 25882 13101 25899
rect 13072 25879 13101 25882
rect 21237 25899 21266 25902
rect 21237 25882 21243 25899
rect 21260 25898 21266 25899
rect 21544 25898 21558 25918
rect 21636 25902 21650 25918
rect 21260 25884 21558 25898
rect 21628 25899 21657 25902
rect 21260 25882 21266 25884
rect 21237 25879 21266 25882
rect 21628 25882 21634 25899
rect 21651 25898 21657 25899
rect 22869 25898 22872 25904
rect 21651 25884 22872 25898
rect 21651 25882 21657 25884
rect 21628 25879 21657 25882
rect 22869 25878 22872 25884
rect 22898 25878 22901 25904
rect 3036 25816 29992 25864
rect 7045 25776 7048 25802
rect 7074 25796 7077 25802
rect 7551 25796 7554 25802
rect 7074 25782 7554 25796
rect 7074 25776 7077 25782
rect 7551 25776 7554 25782
rect 7580 25796 7583 25802
rect 9070 25797 9099 25800
rect 7580 25782 9046 25796
rect 7580 25776 7583 25782
rect 8978 25763 9007 25766
rect 8978 25746 8984 25763
rect 9001 25746 9007 25763
rect 9032 25762 9046 25782
rect 9070 25780 9076 25797
rect 9093 25796 9099 25797
rect 9253 25796 9256 25802
rect 9093 25782 9256 25796
rect 9093 25780 9099 25782
rect 9070 25777 9099 25780
rect 9253 25776 9256 25782
rect 9282 25776 9285 25802
rect 16291 25776 16294 25802
rect 16320 25796 16323 25802
rect 16384 25797 16413 25800
rect 16384 25796 16390 25797
rect 16320 25782 16390 25796
rect 16320 25776 16323 25782
rect 16384 25780 16390 25782
rect 16407 25780 16413 25797
rect 16384 25777 16413 25780
rect 17487 25776 17490 25802
rect 17516 25776 17519 25802
rect 23007 25776 23010 25802
rect 23036 25776 23039 25802
rect 9032 25748 9184 25762
rect 8978 25743 9007 25746
rect 7229 25708 7232 25734
rect 7258 25728 7261 25734
rect 8986 25728 9000 25743
rect 9170 25732 9184 25748
rect 7258 25714 7850 25728
rect 7258 25708 7261 25714
rect 4654 25695 4683 25698
rect 4654 25678 4660 25695
rect 4677 25694 4683 25695
rect 4699 25694 4702 25700
rect 4677 25680 4702 25694
rect 4677 25678 4683 25680
rect 4654 25675 4683 25678
rect 4699 25674 4702 25680
rect 4728 25674 4731 25700
rect 4791 25674 4794 25700
rect 4820 25698 4823 25700
rect 4820 25695 4838 25698
rect 4832 25678 4838 25695
rect 4820 25675 4838 25678
rect 4853 25695 4882 25698
rect 4853 25678 4859 25695
rect 4876 25694 4882 25695
rect 5205 25694 5208 25700
rect 4876 25680 5208 25694
rect 4876 25678 4882 25680
rect 4853 25675 4882 25678
rect 4820 25674 4823 25675
rect 5205 25674 5208 25680
rect 5234 25674 5237 25700
rect 7735 25674 7738 25700
rect 7764 25674 7767 25700
rect 7836 25698 7850 25714
rect 8250 25714 9000 25728
rect 9162 25729 9191 25732
rect 8250 25698 8264 25714
rect 9162 25712 9168 25729
rect 9185 25712 9191 25729
rect 9162 25709 9191 25712
rect 13716 25729 13745 25732
rect 13716 25712 13722 25729
rect 13739 25728 13745 25729
rect 16154 25729 16183 25732
rect 16154 25728 16160 25729
rect 13739 25714 16160 25728
rect 13739 25712 13745 25714
rect 13716 25709 13745 25712
rect 16154 25712 16160 25714
rect 16177 25712 16183 25729
rect 16154 25709 16183 25712
rect 17119 25708 17122 25734
rect 17148 25728 17151 25734
rect 17258 25729 17287 25732
rect 17258 25728 17264 25729
rect 17148 25714 17264 25728
rect 17148 25708 17151 25714
rect 17258 25712 17264 25714
rect 17281 25712 17287 25729
rect 17258 25709 17287 25712
rect 23054 25729 23083 25732
rect 23054 25712 23060 25729
rect 23077 25728 23083 25729
rect 23651 25728 23654 25734
rect 23077 25714 23654 25728
rect 23077 25712 23083 25714
rect 23054 25709 23083 25712
rect 23651 25708 23654 25714
rect 23680 25708 23683 25734
rect 7828 25695 7857 25698
rect 7828 25678 7834 25695
rect 7851 25678 7857 25695
rect 7828 25675 7857 25678
rect 8242 25695 8271 25698
rect 8242 25678 8248 25695
rect 8265 25678 8271 25695
rect 8242 25675 8271 25678
rect 8334 25695 8363 25698
rect 8334 25678 8340 25695
rect 8357 25678 8363 25695
rect 8334 25675 8363 25678
rect 7782 25661 7811 25664
rect 7782 25644 7788 25661
rect 7805 25660 7811 25661
rect 8342 25660 8356 25675
rect 8517 25674 8520 25700
rect 8546 25674 8549 25700
rect 8748 25695 8777 25698
rect 8748 25678 8754 25695
rect 8771 25694 8777 25695
rect 8771 25680 9092 25694
rect 8771 25678 8777 25680
rect 8748 25675 8777 25678
rect 7805 25646 8356 25660
rect 8978 25661 9007 25664
rect 7805 25644 7811 25646
rect 7782 25641 7811 25644
rect 8978 25644 8984 25661
rect 9001 25644 9007 25661
rect 8978 25641 9007 25644
rect 5689 25627 5718 25630
rect 5689 25610 5695 25627
rect 5712 25626 5718 25627
rect 6171 25626 6174 25632
rect 5712 25612 6174 25626
rect 5712 25610 5718 25612
rect 5689 25607 5718 25610
rect 6171 25606 6174 25612
rect 6200 25606 6203 25632
rect 8103 25606 8106 25632
rect 8132 25626 8135 25632
rect 8241 25626 8244 25632
rect 8132 25612 8244 25626
rect 8132 25606 8135 25612
rect 8241 25606 8244 25612
rect 8270 25626 8273 25632
rect 8986 25626 9000 25641
rect 8270 25612 9000 25626
rect 9078 25626 9092 25680
rect 9115 25674 9118 25700
rect 9144 25694 9147 25700
rect 9575 25694 9578 25700
rect 9144 25680 9578 25694
rect 9144 25674 9147 25680
rect 9575 25674 9578 25680
rect 9604 25674 9607 25700
rect 12979 25674 12982 25700
rect 13008 25694 13011 25700
rect 13485 25694 13488 25700
rect 13008 25680 13488 25694
rect 13008 25674 13011 25680
rect 13485 25674 13488 25680
rect 13514 25694 13517 25700
rect 13670 25695 13699 25698
rect 13670 25694 13676 25695
rect 13514 25680 13676 25694
rect 13514 25674 13517 25680
rect 13670 25678 13676 25680
rect 13693 25678 13699 25695
rect 13670 25675 13699 25678
rect 13762 25695 13791 25698
rect 13762 25678 13768 25695
rect 13785 25678 13791 25695
rect 13762 25675 13791 25678
rect 16200 25695 16229 25698
rect 16200 25678 16206 25695
rect 16223 25678 16229 25695
rect 16200 25675 16229 25678
rect 13531 25640 13534 25666
rect 13560 25660 13563 25666
rect 13770 25660 13784 25675
rect 13560 25646 13784 25660
rect 16208 25660 16222 25675
rect 16705 25674 16708 25700
rect 16734 25694 16737 25700
rect 17211 25694 17214 25700
rect 16734 25680 17214 25694
rect 16734 25674 16737 25680
rect 17211 25674 17214 25680
rect 17240 25694 17243 25700
rect 17304 25695 17333 25698
rect 17304 25694 17310 25695
rect 17240 25680 17310 25694
rect 17240 25674 17243 25680
rect 17304 25678 17310 25680
rect 17327 25678 17333 25695
rect 17304 25675 17333 25678
rect 20477 25674 20480 25700
rect 20506 25694 20509 25700
rect 20570 25695 20599 25698
rect 20570 25694 20576 25695
rect 20506 25680 20576 25694
rect 20506 25674 20509 25680
rect 20570 25678 20576 25680
rect 20593 25678 20599 25695
rect 20570 25675 20599 25678
rect 21535 25674 21538 25700
rect 21564 25694 21567 25700
rect 21582 25695 21611 25698
rect 21582 25694 21588 25695
rect 21564 25680 21588 25694
rect 21564 25674 21567 25680
rect 21582 25678 21588 25680
rect 21605 25678 21611 25695
rect 22824 25695 22853 25698
rect 22824 25694 22830 25695
rect 21582 25675 21611 25678
rect 22763 25680 22830 25694
rect 17257 25660 17260 25666
rect 16208 25646 17260 25660
rect 13560 25640 13563 25646
rect 17257 25640 17260 25646
rect 17286 25640 17289 25666
rect 22763 25660 22777 25680
rect 22824 25678 22830 25680
rect 22847 25678 22853 25695
rect 22824 25675 22853 25678
rect 22869 25674 22872 25700
rect 22898 25674 22901 25700
rect 23099 25674 23102 25700
rect 23128 25674 23131 25700
rect 21360 25646 22777 25660
rect 21360 25632 21374 25646
rect 15923 25626 15926 25632
rect 9078 25612 15926 25626
rect 8270 25606 8273 25612
rect 15923 25606 15926 25612
rect 15952 25606 15955 25632
rect 20616 25627 20645 25630
rect 20616 25610 20622 25627
rect 20639 25626 20645 25627
rect 21351 25626 21354 25632
rect 20639 25612 21354 25626
rect 20639 25610 20645 25612
rect 20616 25607 20645 25610
rect 21351 25606 21354 25612
rect 21380 25606 21383 25632
rect 21443 25606 21446 25632
rect 21472 25626 21475 25632
rect 21581 25626 21584 25632
rect 21472 25612 21584 25626
rect 21472 25606 21475 25612
rect 21581 25606 21584 25612
rect 21610 25626 21613 25632
rect 21628 25627 21657 25630
rect 21628 25626 21634 25627
rect 21610 25612 21634 25626
rect 21610 25606 21613 25612
rect 21628 25610 21634 25612
rect 21651 25610 21657 25627
rect 21628 25607 21657 25610
rect 3036 25544 29992 25592
rect 4883 25504 4886 25530
rect 4912 25524 4915 25530
rect 5527 25524 5530 25530
rect 4912 25510 5530 25524
rect 4912 25504 4915 25510
rect 5527 25504 5530 25510
rect 5556 25504 5559 25530
rect 7551 25528 7554 25530
rect 7529 25525 7554 25528
rect 7529 25508 7535 25525
rect 7552 25508 7554 25525
rect 7529 25505 7554 25508
rect 7551 25504 7554 25505
rect 7580 25504 7583 25530
rect 8058 25525 8087 25528
rect 8058 25508 8064 25525
rect 8081 25524 8087 25525
rect 8517 25524 8520 25530
rect 8081 25510 8520 25524
rect 8081 25508 8087 25510
rect 8058 25505 8087 25508
rect 8517 25504 8520 25510
rect 8546 25504 8549 25530
rect 8655 25504 8658 25530
rect 8684 25524 8687 25530
rect 8839 25524 8842 25530
rect 8684 25510 8842 25524
rect 8684 25504 8687 25510
rect 8839 25504 8842 25510
rect 8868 25524 8871 25530
rect 9621 25524 9624 25530
rect 8868 25510 9624 25524
rect 8868 25504 8871 25510
rect 9621 25504 9624 25510
rect 9650 25504 9653 25530
rect 18867 25504 18870 25530
rect 18896 25504 18899 25530
rect 23651 25504 23654 25530
rect 23680 25504 23683 25530
rect 3273 25470 3276 25496
rect 3302 25490 3305 25496
rect 6705 25491 6734 25494
rect 3302 25476 3480 25490
rect 3302 25470 3305 25476
rect 3366 25457 3395 25460
rect 3366 25440 3372 25457
rect 3389 25456 3395 25457
rect 3411 25456 3414 25462
rect 3389 25442 3414 25456
rect 3389 25440 3395 25442
rect 3366 25437 3395 25440
rect 3411 25436 3414 25442
rect 3440 25436 3443 25462
rect 3466 25456 3480 25476
rect 6705 25474 6711 25491
rect 6728 25490 6734 25491
rect 6769 25490 6772 25496
rect 6728 25476 6772 25490
rect 6728 25474 6734 25476
rect 6705 25471 6734 25474
rect 6769 25470 6772 25476
rect 6798 25470 6801 25496
rect 9032 25476 9888 25490
rect 3521 25457 3550 25460
rect 3521 25456 3527 25457
rect 3466 25442 3527 25456
rect 3521 25440 3527 25442
rect 3544 25440 3550 25457
rect 3521 25437 3550 25440
rect 3565 25457 3594 25460
rect 3565 25440 3571 25457
rect 3588 25456 3594 25457
rect 3641 25456 3644 25462
rect 3588 25442 3644 25456
rect 3588 25440 3594 25442
rect 3565 25437 3594 25440
rect 3641 25436 3644 25442
rect 3670 25436 3673 25462
rect 5527 25436 5530 25462
rect 5556 25456 5559 25462
rect 6494 25457 6523 25460
rect 6494 25456 6500 25457
rect 5556 25442 6500 25456
rect 5556 25436 5559 25442
rect 6494 25440 6500 25442
rect 6517 25440 6523 25457
rect 6494 25437 6523 25440
rect 6631 25436 6634 25462
rect 6660 25460 6663 25462
rect 6660 25457 6678 25460
rect 6672 25440 6678 25457
rect 8058 25457 8087 25460
rect 8058 25456 8064 25457
rect 6660 25437 6678 25440
rect 7422 25442 8064 25456
rect 6660 25436 6663 25437
rect 7422 25428 7436 25442
rect 8058 25440 8064 25442
rect 8081 25440 8087 25457
rect 8058 25437 8087 25440
rect 7413 25402 7416 25428
rect 7442 25402 7445 25428
rect 8196 25423 8225 25426
rect 8196 25406 8202 25423
rect 8219 25422 8225 25423
rect 8333 25422 8336 25428
rect 8219 25408 8336 25422
rect 8219 25406 8225 25408
rect 8196 25403 8225 25406
rect 8333 25402 8336 25408
rect 8362 25422 8365 25428
rect 8931 25422 8934 25428
rect 8362 25408 8934 25422
rect 8362 25402 8365 25408
rect 8931 25402 8934 25408
rect 8960 25402 8963 25428
rect 4469 25368 4472 25394
rect 4498 25388 4501 25394
rect 4498 25374 6217 25388
rect 4498 25368 4501 25374
rect 4401 25355 4430 25358
rect 4401 25338 4407 25355
rect 4424 25354 4430 25355
rect 4791 25354 4794 25360
rect 4424 25340 4794 25354
rect 4424 25338 4430 25340
rect 4401 25335 4430 25338
rect 4791 25334 4794 25340
rect 4820 25334 4823 25360
rect 6203 25354 6217 25374
rect 8057 25368 8060 25394
rect 8086 25388 8089 25394
rect 8104 25389 8133 25392
rect 8104 25388 8110 25389
rect 8086 25374 8110 25388
rect 8086 25368 8089 25374
rect 8104 25372 8110 25374
rect 8127 25388 8133 25389
rect 8149 25388 8152 25394
rect 8127 25374 8152 25388
rect 8127 25372 8133 25374
rect 8104 25369 8133 25372
rect 8149 25368 8152 25374
rect 8178 25368 8181 25394
rect 9032 25354 9046 25476
rect 9069 25436 9072 25462
rect 9098 25456 9101 25462
rect 9874 25460 9888 25476
rect 18315 25470 18318 25496
rect 18344 25490 18347 25496
rect 19190 25491 19219 25494
rect 19190 25490 19196 25491
rect 18344 25476 19196 25490
rect 18344 25470 18347 25476
rect 19190 25474 19196 25476
rect 19213 25474 19219 25491
rect 19190 25471 19219 25474
rect 9823 25457 9852 25460
rect 9823 25456 9829 25457
rect 9098 25442 9829 25456
rect 9098 25436 9101 25442
rect 9823 25440 9829 25442
rect 9846 25440 9852 25457
rect 9823 25437 9852 25440
rect 9867 25457 9896 25460
rect 9867 25440 9873 25457
rect 9890 25456 9896 25457
rect 10679 25456 10682 25462
rect 9890 25442 10682 25456
rect 9890 25440 9896 25442
rect 9867 25437 9896 25440
rect 10679 25436 10682 25442
rect 10708 25436 10711 25462
rect 17901 25436 17904 25462
rect 17930 25456 17933 25462
rect 18684 25457 18713 25460
rect 18684 25456 18690 25457
rect 17930 25442 18690 25456
rect 17930 25436 17933 25442
rect 18684 25440 18690 25442
rect 18707 25440 18713 25457
rect 18684 25437 18713 25440
rect 18775 25436 18778 25462
rect 18804 25456 18807 25462
rect 19098 25457 19127 25460
rect 19098 25456 19104 25457
rect 18804 25442 19104 25456
rect 18804 25436 18807 25442
rect 19098 25440 19104 25442
rect 19121 25440 19127 25457
rect 19098 25437 19127 25440
rect 19236 25457 19265 25460
rect 19236 25440 19242 25457
rect 19259 25440 19265 25457
rect 19236 25437 19265 25440
rect 9668 25423 9697 25426
rect 9668 25406 9674 25423
rect 9691 25406 9697 25423
rect 9668 25403 9697 25406
rect 18730 25423 18759 25426
rect 18730 25406 18736 25423
rect 18753 25422 18759 25423
rect 18913 25422 18916 25428
rect 18753 25408 18916 25422
rect 18753 25406 18759 25408
rect 18730 25403 18759 25406
rect 6203 25340 9046 25354
rect 9621 25334 9624 25360
rect 9650 25354 9653 25360
rect 9676 25354 9690 25403
rect 18913 25402 18916 25408
rect 18942 25422 18945 25428
rect 19244 25422 19258 25437
rect 23329 25436 23332 25462
rect 23358 25456 23361 25462
rect 23514 25457 23543 25460
rect 23514 25456 23520 25457
rect 23358 25442 23520 25456
rect 23358 25436 23361 25442
rect 23514 25440 23520 25442
rect 23537 25440 23543 25457
rect 23514 25437 23543 25440
rect 18942 25408 19258 25422
rect 18942 25402 18945 25408
rect 23283 25402 23286 25428
rect 23312 25422 23315 25428
rect 23422 25423 23451 25426
rect 23422 25422 23428 25423
rect 23312 25408 23428 25422
rect 23312 25402 23315 25408
rect 23422 25406 23428 25408
rect 23445 25406 23451 25423
rect 23422 25403 23451 25406
rect 23698 25423 23727 25426
rect 23698 25406 23704 25423
rect 23721 25406 23727 25423
rect 23698 25403 23727 25406
rect 11047 25388 11050 25394
rect 10504 25374 11050 25388
rect 10504 25354 10518 25374
rect 11047 25368 11050 25374
rect 11076 25368 11079 25394
rect 23099 25368 23102 25394
rect 23128 25388 23131 25394
rect 23706 25388 23720 25403
rect 23128 25374 23720 25388
rect 23128 25368 23131 25374
rect 9650 25340 10518 25354
rect 10703 25355 10732 25358
rect 9650 25334 9653 25340
rect 10703 25338 10709 25355
rect 10726 25354 10732 25355
rect 10771 25354 10774 25360
rect 10726 25340 10774 25354
rect 10726 25338 10732 25340
rect 10703 25335 10732 25338
rect 10771 25334 10774 25340
rect 10800 25334 10803 25360
rect 19097 25334 19100 25360
rect 19126 25334 19129 25360
rect 23559 25334 23562 25360
rect 23588 25334 23591 25360
rect 3036 25272 29992 25320
rect 3411 25252 3414 25258
rect 3144 25238 3414 25252
rect 3144 25188 3158 25238
rect 3411 25232 3414 25238
rect 3440 25232 3443 25258
rect 8149 25232 8152 25258
rect 8178 25252 8181 25258
rect 8178 25238 9552 25252
rect 8178 25232 8181 25238
rect 3136 25185 3165 25188
rect 3136 25168 3142 25185
rect 3159 25168 3165 25185
rect 9538 25184 9552 25238
rect 11231 25232 11234 25258
rect 11260 25252 11263 25258
rect 12841 25252 12844 25258
rect 11260 25238 12844 25252
rect 11260 25232 11263 25238
rect 12841 25232 12844 25238
rect 12870 25232 12873 25258
rect 17395 25232 17398 25258
rect 17424 25232 17427 25258
rect 22709 25253 22738 25256
rect 22709 25236 22715 25253
rect 22732 25252 22738 25253
rect 23099 25252 23102 25258
rect 22732 25238 23102 25252
rect 22732 25236 22738 25238
rect 22709 25233 22738 25236
rect 23099 25232 23102 25238
rect 23128 25232 23131 25258
rect 15049 25184 15052 25190
rect 3136 25165 3165 25168
rect 4110 25170 8724 25184
rect 9538 25170 11070 25184
rect 3273 25130 3276 25156
rect 3302 25154 3305 25156
rect 3302 25151 3320 25154
rect 3314 25134 3320 25151
rect 3733 25150 3736 25156
rect 3302 25131 3320 25134
rect 3466 25136 3736 25150
rect 3302 25130 3305 25131
rect 3347 25117 3376 25120
rect 3347 25100 3353 25117
rect 3370 25116 3376 25117
rect 3466 25116 3480 25136
rect 3733 25130 3736 25136
rect 3762 25150 3765 25156
rect 4110 25150 4124 25170
rect 3762 25136 4124 25150
rect 4171 25151 4200 25154
rect 3762 25130 3765 25136
rect 4171 25134 4177 25151
rect 4194 25150 4200 25151
rect 4654 25151 4683 25154
rect 4654 25150 4660 25151
rect 4194 25136 4660 25150
rect 4194 25134 4200 25136
rect 4171 25131 4200 25134
rect 4654 25134 4660 25136
rect 4677 25134 4683 25151
rect 4654 25131 4683 25134
rect 4791 25130 4794 25156
rect 4820 25130 4823 25156
rect 4838 25151 4867 25154
rect 4838 25134 4844 25151
rect 4861 25150 4867 25151
rect 5251 25150 5254 25156
rect 4861 25136 5254 25150
rect 4861 25134 4867 25136
rect 4838 25131 4867 25134
rect 5251 25130 5254 25136
rect 5280 25130 5283 25156
rect 8287 25130 8290 25156
rect 8316 25150 8319 25156
rect 8655 25150 8658 25156
rect 8316 25136 8658 25150
rect 8316 25130 8319 25136
rect 8655 25130 8658 25136
rect 8684 25130 8687 25156
rect 8710 25150 8724 25170
rect 8710 25136 9690 25150
rect 3370 25102 3480 25116
rect 4746 25117 4775 25120
rect 3370 25100 3376 25102
rect 3347 25097 3376 25100
rect 4746 25100 4752 25117
rect 4769 25116 4775 25117
rect 4883 25116 4886 25122
rect 4769 25102 4886 25116
rect 4769 25100 4775 25102
rect 4746 25097 4775 25100
rect 4883 25096 4886 25102
rect 4912 25096 4915 25122
rect 8333 25096 8336 25122
rect 8362 25116 8365 25122
rect 8894 25120 8908 25136
rect 8816 25117 8845 25120
rect 8816 25116 8822 25117
rect 8362 25102 8822 25116
rect 8362 25096 8365 25102
rect 8816 25100 8822 25102
rect 8839 25100 8845 25117
rect 8816 25097 8845 25100
rect 8867 25117 8908 25120
rect 8867 25100 8873 25117
rect 8890 25102 8908 25117
rect 9676 25116 9690 25136
rect 11001 25130 11004 25156
rect 11030 25130 11033 25156
rect 11056 25150 11070 25170
rect 14874 25170 15052 25184
rect 11163 25151 11192 25154
rect 11163 25150 11169 25151
rect 11056 25136 11169 25150
rect 11163 25134 11169 25136
rect 11186 25150 11192 25151
rect 11323 25150 11326 25156
rect 11186 25136 11326 25150
rect 11186 25134 11192 25136
rect 11163 25131 11192 25134
rect 11323 25130 11326 25136
rect 11352 25130 11355 25156
rect 14874 25154 14888 25170
rect 15049 25164 15052 25170
rect 15078 25164 15081 25190
rect 17073 25164 17076 25190
rect 17102 25184 17105 25190
rect 17166 25185 17195 25188
rect 17166 25184 17172 25185
rect 17102 25170 17172 25184
rect 17102 25164 17105 25170
rect 17166 25168 17172 25170
rect 17189 25168 17195 25185
rect 17166 25165 17195 25168
rect 18361 25164 18364 25190
rect 18390 25184 18393 25190
rect 18499 25184 18502 25190
rect 18390 25170 18502 25184
rect 18390 25164 18393 25170
rect 18499 25164 18502 25170
rect 18528 25164 18531 25190
rect 20386 25185 20415 25188
rect 20386 25168 20392 25185
rect 20409 25184 20415 25185
rect 20409 25170 21742 25184
rect 20409 25168 20415 25170
rect 20386 25165 20415 25168
rect 14866 25151 14895 25154
rect 14866 25134 14872 25151
rect 14889 25134 14895 25151
rect 14866 25131 14895 25134
rect 14911 25130 14914 25156
rect 14940 25130 14943 25156
rect 14958 25151 14987 25154
rect 14958 25134 14964 25151
rect 14981 25150 14987 25151
rect 15003 25150 15006 25156
rect 14981 25136 15006 25150
rect 14981 25134 14987 25136
rect 14958 25131 14987 25134
rect 15003 25130 15006 25136
rect 15032 25130 15035 25156
rect 16153 25130 16156 25156
rect 16182 25150 16185 25156
rect 17212 25151 17241 25154
rect 17212 25150 17218 25151
rect 16182 25136 17218 25150
rect 16182 25130 16185 25136
rect 11231 25120 11234 25122
rect 11213 25117 11234 25120
rect 11213 25116 11219 25117
rect 9676 25102 11219 25116
rect 8890 25100 8896 25102
rect 8867 25097 8896 25100
rect 11213 25100 11219 25102
rect 11213 25097 11234 25100
rect 11231 25096 11234 25097
rect 11260 25096 11263 25122
rect 4930 25083 4959 25086
rect 4930 25066 4936 25083
rect 4953 25082 4959 25083
rect 6355 25082 6358 25088
rect 4953 25068 6358 25082
rect 4953 25066 4959 25068
rect 4930 25063 4959 25066
rect 6355 25062 6358 25068
rect 6384 25062 6387 25088
rect 9691 25083 9720 25086
rect 9691 25066 9697 25083
rect 9714 25082 9720 25083
rect 10495 25082 10498 25088
rect 9714 25068 10498 25082
rect 9714 25066 9720 25068
rect 9691 25063 9720 25066
rect 10495 25062 10498 25068
rect 10524 25062 10527 25088
rect 12059 25086 12062 25088
rect 12037 25083 12062 25086
rect 12037 25066 12043 25083
rect 12060 25066 12062 25083
rect 12037 25063 12062 25066
rect 12059 25062 12062 25063
rect 12088 25062 12091 25088
rect 14497 25062 14500 25088
rect 14526 25082 14529 25088
rect 15050 25083 15079 25086
rect 15050 25082 15056 25083
rect 14526 25068 15056 25082
rect 14526 25062 14529 25068
rect 15050 25066 15056 25068
rect 15073 25066 15079 25083
rect 17128 25082 17142 25136
rect 17212 25134 17218 25136
rect 17235 25134 17241 25151
rect 17764 25151 17793 25154
rect 17764 25150 17770 25151
rect 17212 25131 17241 25134
rect 17266 25136 17770 25150
rect 17165 25096 17168 25122
rect 17194 25116 17197 25122
rect 17266 25116 17280 25136
rect 17764 25134 17770 25136
rect 17787 25134 17793 25151
rect 17764 25131 17793 25134
rect 18634 25151 18663 25154
rect 18634 25134 18640 25151
rect 18657 25150 18663 25151
rect 19097 25150 19100 25156
rect 18657 25136 19100 25150
rect 18657 25134 18663 25136
rect 18634 25131 18663 25134
rect 19097 25130 19100 25136
rect 19126 25130 19129 25156
rect 20340 25151 20369 25154
rect 20340 25134 20346 25151
rect 20363 25150 20369 25151
rect 20477 25150 20480 25156
rect 20363 25136 20480 25150
rect 20363 25134 20369 25136
rect 20340 25131 20369 25134
rect 20477 25130 20480 25136
rect 20506 25130 20509 25156
rect 21673 25130 21676 25156
rect 21702 25130 21705 25156
rect 21728 25150 21742 25170
rect 21835 25151 21864 25154
rect 21835 25150 21841 25151
rect 21728 25136 21841 25150
rect 21835 25134 21841 25136
rect 21858 25150 21864 25151
rect 23927 25150 23930 25156
rect 21858 25136 23930 25150
rect 21858 25134 21864 25136
rect 21835 25131 21864 25134
rect 23927 25130 23930 25136
rect 23956 25130 23959 25156
rect 17194 25102 17280 25116
rect 17626 25117 17655 25120
rect 17194 25096 17197 25102
rect 17626 25100 17632 25117
rect 17649 25100 17655 25117
rect 17626 25097 17655 25100
rect 17634 25082 17648 25097
rect 17717 25096 17720 25122
rect 17746 25096 17749 25122
rect 18545 25096 18548 25122
rect 18574 25116 18577 25122
rect 21903 25120 21906 25122
rect 21885 25117 21906 25120
rect 18574 25102 19212 25116
rect 18574 25096 18577 25102
rect 17128 25068 17648 25082
rect 17764 25083 17793 25086
rect 15050 25063 15079 25066
rect 17764 25066 17770 25083
rect 17787 25082 17793 25083
rect 18683 25082 18686 25088
rect 17787 25068 18686 25082
rect 17787 25066 17793 25068
rect 17764 25063 17793 25066
rect 18683 25062 18686 25068
rect 18712 25062 18715 25088
rect 19198 25086 19212 25102
rect 21885 25100 21891 25117
rect 21885 25097 21906 25100
rect 21903 25096 21906 25097
rect 21932 25096 21935 25122
rect 19190 25083 19219 25086
rect 19190 25066 19196 25083
rect 19213 25066 19219 25083
rect 19190 25063 19219 25066
rect 20385 25062 20388 25088
rect 20414 25082 20417 25088
rect 20524 25083 20553 25086
rect 20524 25082 20530 25083
rect 20414 25068 20530 25082
rect 20414 25062 20417 25068
rect 20524 25066 20530 25068
rect 20547 25066 20553 25083
rect 20524 25063 20553 25066
rect 3036 25000 29992 25048
rect 12888 24981 12917 24984
rect 12888 24964 12894 24981
rect 12911 24964 12917 24981
rect 15003 24980 15006 24986
rect 12888 24961 12917 24964
rect 14874 24966 15006 24980
rect 9667 24926 9670 24952
rect 9696 24946 9699 24952
rect 9821 24947 9850 24950
rect 9821 24946 9827 24947
rect 9696 24932 9827 24946
rect 9696 24926 9699 24932
rect 9821 24930 9827 24932
rect 9844 24930 9850 24947
rect 9821 24927 9850 24930
rect 10679 24926 10682 24952
rect 10708 24946 10711 24952
rect 11765 24947 11794 24950
rect 11765 24946 11771 24947
rect 10708 24932 11771 24946
rect 10708 24926 10711 24932
rect 11765 24930 11771 24932
rect 11788 24946 11794 24947
rect 11788 24930 11806 24946
rect 11765 24927 11806 24930
rect 5803 24892 5806 24918
rect 5832 24912 5835 24918
rect 6034 24913 6063 24916
rect 6034 24912 6040 24913
rect 5832 24898 6040 24912
rect 5832 24892 5835 24898
rect 6034 24896 6040 24898
rect 6057 24896 6063 24913
rect 6034 24893 6063 24896
rect 6079 24892 6082 24918
rect 6108 24916 6111 24918
rect 6108 24913 6120 24916
rect 6114 24896 6120 24913
rect 6108 24893 6120 24896
rect 6108 24892 6111 24893
rect 6171 24892 6174 24918
rect 6200 24916 6203 24918
rect 6200 24913 6214 24916
rect 6208 24896 6214 24913
rect 6295 24913 6324 24916
rect 6200 24893 6214 24896
rect 6240 24908 6269 24911
rect 6200 24892 6203 24893
rect 6240 24891 6246 24908
rect 6263 24891 6269 24908
rect 6295 24896 6301 24913
rect 6318 24912 6324 24913
rect 6346 24913 6375 24916
rect 6318 24896 6332 24912
rect 6295 24893 6332 24896
rect 6346 24896 6352 24913
rect 6369 24912 6375 24913
rect 7781 24912 7784 24918
rect 6369 24898 7784 24912
rect 6369 24896 6375 24898
rect 6346 24893 6375 24896
rect 6240 24888 6269 24891
rect 6248 24844 6262 24888
rect 6318 24878 6332 24893
rect 7781 24892 7784 24898
rect 7810 24892 7813 24918
rect 8931 24892 8934 24918
rect 8960 24912 8963 24918
rect 9777 24913 9806 24916
rect 9777 24912 9783 24913
rect 8960 24898 9783 24912
rect 8960 24892 8963 24898
rect 9777 24896 9783 24898
rect 9800 24896 9806 24913
rect 9777 24893 9806 24896
rect 11369 24892 11372 24918
rect 11398 24912 11401 24918
rect 11709 24913 11738 24916
rect 11709 24912 11715 24913
rect 11398 24898 11715 24912
rect 11398 24892 11401 24898
rect 11709 24896 11715 24898
rect 11732 24896 11738 24913
rect 11792 24912 11806 24927
rect 12795 24912 12798 24918
rect 11792 24898 12798 24912
rect 11709 24893 11738 24896
rect 12795 24892 12798 24898
rect 12824 24892 12827 24918
rect 6539 24878 6542 24884
rect 6318 24864 6542 24878
rect 6539 24858 6542 24864
rect 6568 24858 6571 24884
rect 9621 24858 9624 24884
rect 9650 24858 9653 24884
rect 11047 24858 11050 24884
rect 11076 24878 11079 24884
rect 11554 24879 11583 24882
rect 11554 24878 11560 24879
rect 11076 24864 11560 24878
rect 11076 24858 11079 24864
rect 11554 24862 11560 24864
rect 11577 24862 11583 24879
rect 11554 24859 11583 24862
rect 6493 24844 6496 24850
rect 6248 24830 6496 24844
rect 6493 24824 6496 24830
rect 6522 24824 6525 24850
rect 12896 24844 12910 24961
rect 12980 24913 13009 24916
rect 12980 24896 12986 24913
rect 13003 24896 13009 24913
rect 12980 24893 13009 24896
rect 12988 24878 13002 24893
rect 13117 24892 13120 24918
rect 13146 24892 13149 24918
rect 13255 24892 13258 24918
rect 13284 24892 13287 24918
rect 13348 24913 13377 24916
rect 13348 24896 13354 24913
rect 13371 24912 13377 24913
rect 13991 24912 13994 24918
rect 13371 24898 13994 24912
rect 13371 24896 13377 24898
rect 13348 24893 13377 24896
rect 13991 24892 13994 24898
rect 14020 24892 14023 24918
rect 14773 24892 14776 24918
rect 14802 24912 14805 24918
rect 14874 24916 14888 24966
rect 15003 24960 15006 24966
rect 15032 24980 15035 24986
rect 15877 24980 15880 24986
rect 15032 24966 15880 24980
rect 15032 24960 15035 24966
rect 15877 24960 15880 24966
rect 15906 24980 15909 24986
rect 18315 24980 18318 24986
rect 15906 24966 18318 24980
rect 15906 24960 15909 24966
rect 18315 24960 18318 24966
rect 18344 24960 18347 24986
rect 14911 24926 14914 24952
rect 14940 24946 14943 24952
rect 14940 24932 15210 24946
rect 14940 24926 14943 24932
rect 15196 24916 15210 24932
rect 15242 24932 18292 24946
rect 14866 24913 14895 24916
rect 14866 24912 14872 24913
rect 14802 24898 14872 24912
rect 14802 24892 14805 24898
rect 14866 24896 14872 24898
rect 14889 24896 14895 24913
rect 14866 24893 14895 24896
rect 15142 24913 15171 24916
rect 15142 24896 15148 24913
rect 15165 24896 15171 24913
rect 15142 24893 15171 24896
rect 15188 24913 15217 24916
rect 15188 24896 15194 24913
rect 15211 24896 15217 24913
rect 15188 24893 15217 24896
rect 12988 24864 13416 24878
rect 12390 24830 12910 24844
rect 13402 24844 13416 24864
rect 15049 24858 15052 24884
rect 15078 24878 15081 24884
rect 15150 24878 15164 24893
rect 15242 24878 15256 24932
rect 15326 24913 15355 24916
rect 15326 24896 15332 24913
rect 15349 24912 15355 24913
rect 15832 24913 15861 24916
rect 15832 24912 15838 24913
rect 15349 24898 15838 24912
rect 15349 24896 15355 24898
rect 15326 24893 15355 24896
rect 15832 24896 15838 24898
rect 15855 24896 15861 24913
rect 15832 24893 15861 24896
rect 15078 24864 15256 24878
rect 15840 24878 15854 24893
rect 15877 24892 15880 24918
rect 15906 24892 15909 24918
rect 15932 24916 15946 24932
rect 15924 24913 15953 24916
rect 15924 24896 15930 24913
rect 15947 24896 15953 24913
rect 15924 24893 15953 24896
rect 17073 24892 17076 24918
rect 17102 24892 17105 24918
rect 17257 24892 17260 24918
rect 17286 24912 17289 24918
rect 18278 24916 18292 24932
rect 17350 24913 17379 24916
rect 17350 24912 17356 24913
rect 17286 24898 17356 24912
rect 17286 24892 17289 24898
rect 17350 24896 17356 24898
rect 17373 24896 17379 24913
rect 17350 24893 17379 24896
rect 18270 24913 18299 24916
rect 18270 24896 18276 24913
rect 18293 24912 18299 24913
rect 18545 24912 18548 24918
rect 18293 24898 18548 24912
rect 18293 24896 18299 24898
rect 18270 24893 18299 24896
rect 18545 24892 18548 24898
rect 18574 24912 18577 24918
rect 18730 24913 18759 24916
rect 18730 24912 18736 24913
rect 18574 24898 18736 24912
rect 18574 24892 18577 24898
rect 18730 24896 18736 24898
rect 18753 24896 18759 24913
rect 18730 24893 18759 24896
rect 20340 24913 20369 24916
rect 20340 24896 20346 24913
rect 20363 24912 20369 24913
rect 20363 24898 20707 24912
rect 20363 24896 20369 24898
rect 20340 24893 20369 24896
rect 17165 24878 17168 24884
rect 15840 24864 17168 24878
rect 15078 24858 15081 24864
rect 17165 24858 17168 24864
rect 17194 24858 17197 24884
rect 18315 24858 18318 24884
rect 18344 24858 18347 24884
rect 18408 24879 18437 24882
rect 18408 24862 18414 24879
rect 18431 24878 18437 24879
rect 18453 24878 18456 24884
rect 18431 24864 18456 24878
rect 18431 24862 18437 24864
rect 18408 24859 18437 24862
rect 18453 24858 18456 24864
rect 18482 24858 18485 24884
rect 18683 24858 18686 24884
rect 18712 24858 18715 24884
rect 18913 24858 18916 24884
rect 18942 24858 18945 24884
rect 20385 24858 20388 24884
rect 20414 24858 20417 24884
rect 13807 24844 13810 24850
rect 13402 24830 13810 24844
rect 6034 24811 6063 24814
rect 6034 24794 6040 24811
rect 6057 24810 6063 24811
rect 6401 24810 6404 24816
rect 6057 24796 6404 24810
rect 6057 24794 6063 24796
rect 6034 24791 6063 24794
rect 6401 24790 6404 24796
rect 6430 24790 6433 24816
rect 10633 24790 10636 24816
rect 10662 24814 10665 24816
rect 10662 24811 10686 24814
rect 10662 24794 10663 24811
rect 10680 24794 10686 24811
rect 10662 24791 10686 24794
rect 10662 24790 10665 24791
rect 11323 24790 11326 24816
rect 11352 24810 11355 24816
rect 12390 24810 12404 24830
rect 13807 24824 13810 24830
rect 13836 24824 13839 24850
rect 18362 24845 18391 24848
rect 18362 24828 18368 24845
rect 18385 24844 18391 24845
rect 18775 24844 18778 24850
rect 18385 24830 18778 24844
rect 18385 24828 18391 24830
rect 18362 24825 18391 24828
rect 18775 24824 18778 24830
rect 18804 24824 18807 24850
rect 20693 24844 20707 24898
rect 21397 24892 21400 24918
rect 21426 24892 21429 24918
rect 21444 24879 21473 24882
rect 21444 24862 21450 24879
rect 21467 24878 21473 24879
rect 21535 24878 21538 24884
rect 21467 24864 21538 24878
rect 21467 24862 21473 24864
rect 21444 24859 21473 24862
rect 21535 24858 21538 24864
rect 21564 24858 21567 24884
rect 21582 24845 21611 24848
rect 21582 24844 21588 24845
rect 20693 24830 21588 24844
rect 21582 24828 21588 24830
rect 21605 24828 21611 24845
rect 21582 24825 21611 24828
rect 11352 24796 12404 24810
rect 11352 24790 11355 24796
rect 12427 24790 12430 24816
rect 12456 24810 12459 24816
rect 12589 24811 12618 24814
rect 12589 24810 12595 24811
rect 12456 24796 12595 24810
rect 12456 24790 12459 24796
rect 12589 24794 12595 24796
rect 12612 24794 12618 24811
rect 12589 24791 12618 24794
rect 13394 24811 13423 24814
rect 13394 24794 13400 24811
rect 13417 24810 13423 24811
rect 14405 24810 14408 24816
rect 13417 24796 14408 24810
rect 13417 24794 13423 24796
rect 13394 24791 13423 24794
rect 14405 24790 14408 24796
rect 14434 24790 14437 24816
rect 14865 24790 14868 24816
rect 14894 24790 14897 24816
rect 16015 24790 16018 24816
rect 16044 24790 16047 24816
rect 17119 24790 17122 24816
rect 17148 24790 17151 24816
rect 20339 24790 20342 24816
rect 20368 24810 20371 24816
rect 20478 24811 20507 24814
rect 20478 24810 20484 24811
rect 20368 24796 20484 24810
rect 20368 24790 20371 24796
rect 20478 24794 20484 24796
rect 20501 24794 20507 24811
rect 20478 24791 20507 24794
rect 3036 24728 29992 24776
rect 5803 24688 5806 24714
rect 5832 24708 5835 24714
rect 5832 24694 6516 24708
rect 5832 24688 5835 24694
rect 6502 24674 6516 24694
rect 6539 24688 6542 24714
rect 6568 24712 6571 24714
rect 6568 24709 6592 24712
rect 6568 24692 6569 24709
rect 6586 24692 6592 24709
rect 12335 24708 12338 24714
rect 6568 24689 6592 24692
rect 8204 24694 12338 24708
rect 6568 24688 6571 24689
rect 8204 24674 8218 24694
rect 10725 24674 10728 24680
rect 6502 24660 8218 24674
rect 10711 24654 10728 24674
rect 10754 24654 10757 24680
rect 10771 24654 10774 24680
rect 10800 24654 10803 24680
rect 6953 24620 6956 24646
rect 6982 24640 6985 24646
rect 7736 24641 7765 24644
rect 7736 24640 7742 24641
rect 6982 24626 7742 24640
rect 6982 24620 6985 24626
rect 7736 24624 7742 24626
rect 7759 24624 7765 24641
rect 7736 24621 7765 24624
rect 10711 24616 10725 24654
rect 10780 24616 10794 24654
rect 10703 24613 10732 24616
rect 5159 24586 5162 24612
rect 5188 24606 5191 24612
rect 5527 24606 5530 24612
rect 5188 24592 5530 24606
rect 5188 24586 5191 24592
rect 5527 24586 5530 24592
rect 5556 24586 5559 24612
rect 5665 24586 5668 24612
rect 5694 24610 5697 24612
rect 5694 24607 5712 24610
rect 5706 24590 5712 24607
rect 6217 24606 6220 24612
rect 5694 24587 5712 24590
rect 5858 24592 6220 24606
rect 5694 24586 5697 24587
rect 5739 24573 5768 24576
rect 5739 24556 5745 24573
rect 5762 24572 5768 24573
rect 5858 24572 5872 24592
rect 6217 24586 6220 24592
rect 6246 24586 6249 24612
rect 7919 24586 7922 24612
rect 7948 24610 7951 24612
rect 7948 24606 7952 24610
rect 7948 24592 7970 24606
rect 7948 24587 7952 24592
rect 7948 24586 7951 24587
rect 8195 24586 8198 24612
rect 8224 24586 8227 24612
rect 8241 24586 8244 24612
rect 8270 24606 8273 24612
rect 8395 24607 8424 24610
rect 8395 24606 8401 24607
rect 8270 24592 8401 24606
rect 8270 24586 8273 24592
rect 8395 24590 8401 24592
rect 8418 24606 8424 24607
rect 9207 24606 9210 24612
rect 8418 24592 9210 24606
rect 8418 24590 8424 24592
rect 8395 24587 8424 24590
rect 9207 24586 9210 24592
rect 9236 24586 9239 24612
rect 10495 24586 10498 24612
rect 10524 24586 10527 24612
rect 10541 24586 10544 24612
rect 10570 24610 10573 24612
rect 10570 24607 10582 24610
rect 10576 24590 10582 24607
rect 10570 24587 10582 24590
rect 10570 24586 10573 24587
rect 10633 24586 10636 24612
rect 10662 24608 10665 24612
rect 10662 24605 10676 24608
rect 10670 24588 10676 24605
rect 10703 24596 10709 24613
rect 10726 24596 10732 24613
rect 10703 24593 10732 24596
rect 10757 24613 10794 24616
rect 10757 24596 10763 24613
rect 10780 24597 10794 24613
rect 10826 24610 10840 24694
rect 12335 24688 12338 24694
rect 12364 24688 12367 24714
rect 18223 24688 18226 24714
rect 18252 24708 18255 24714
rect 18684 24709 18713 24712
rect 18684 24708 18690 24709
rect 18252 24694 18690 24708
rect 18252 24688 18255 24694
rect 18684 24692 18690 24694
rect 18707 24692 18713 24709
rect 18684 24689 18713 24692
rect 22985 24709 23014 24712
rect 22985 24692 22991 24709
rect 23008 24708 23014 24709
rect 23329 24708 23332 24714
rect 23008 24694 23332 24708
rect 23008 24692 23014 24694
rect 22985 24689 23014 24692
rect 23329 24688 23332 24694
rect 23358 24688 23361 24714
rect 23651 24688 23654 24714
rect 23680 24708 23683 24714
rect 24020 24709 24049 24712
rect 24020 24708 24026 24709
rect 23680 24694 24026 24708
rect 23680 24688 23683 24694
rect 24020 24692 24026 24694
rect 24043 24692 24049 24709
rect 24020 24689 24049 24692
rect 15832 24675 15861 24678
rect 15832 24674 15838 24675
rect 14483 24660 15838 24674
rect 12381 24620 12384 24646
rect 12410 24640 12413 24646
rect 14483 24640 14497 24660
rect 15832 24658 15838 24660
rect 15855 24658 15861 24675
rect 15832 24655 15861 24658
rect 12410 24626 14497 24640
rect 12410 24620 12413 24626
rect 14773 24620 14776 24646
rect 14802 24620 14805 24646
rect 14911 24620 14914 24646
rect 14940 24640 14943 24646
rect 15004 24641 15033 24644
rect 15004 24640 15010 24641
rect 14940 24626 15010 24640
rect 14940 24620 14943 24626
rect 15004 24624 15010 24626
rect 15027 24624 15033 24641
rect 15004 24621 15033 24624
rect 15049 24620 15052 24646
rect 15078 24620 15081 24646
rect 17257 24640 17260 24646
rect 16944 24626 17260 24640
rect 10808 24607 10840 24610
rect 10780 24596 10786 24597
rect 10757 24593 10786 24596
rect 10662 24586 10676 24588
rect 10808 24590 10814 24607
rect 10831 24592 10840 24607
rect 10831 24590 10837 24592
rect 10808 24587 10837 24590
rect 11047 24586 11050 24612
rect 11076 24606 11079 24612
rect 11094 24607 11123 24610
rect 11094 24606 11100 24607
rect 11076 24592 11100 24606
rect 11076 24586 11079 24592
rect 11094 24590 11100 24592
rect 11117 24590 11123 24607
rect 11094 24587 11123 24590
rect 11255 24607 11284 24610
rect 11255 24590 11261 24607
rect 11278 24606 11284 24607
rect 11369 24606 11372 24612
rect 11278 24592 11372 24606
rect 11278 24590 11284 24592
rect 11255 24587 11284 24590
rect 11369 24586 11372 24592
rect 11398 24586 11401 24612
rect 12979 24586 12982 24612
rect 13008 24606 13011 24612
rect 13026 24607 13055 24610
rect 13026 24606 13032 24607
rect 13008 24592 13032 24606
rect 13008 24586 13011 24592
rect 13026 24590 13032 24592
rect 13049 24590 13055 24607
rect 13026 24587 13055 24590
rect 13302 24607 13331 24610
rect 13302 24590 13308 24607
rect 13325 24590 13331 24607
rect 13302 24587 13331 24590
rect 13762 24607 13791 24610
rect 13762 24590 13768 24607
rect 13785 24606 13791 24607
rect 13807 24606 13810 24612
rect 13785 24592 13810 24606
rect 13785 24590 13791 24592
rect 13762 24587 13791 24590
rect 10647 24585 10676 24586
rect 5762 24558 5872 24572
rect 5762 24556 5768 24558
rect 5739 24553 5768 24556
rect 7735 24552 7738 24578
rect 7764 24552 7767 24578
rect 7828 24573 7857 24576
rect 7828 24556 7834 24573
rect 7851 24556 7857 24573
rect 7828 24553 7857 24556
rect 7836 24538 7850 24553
rect 7873 24552 7876 24578
rect 7902 24552 7905 24578
rect 11323 24576 11326 24578
rect 8356 24573 8385 24576
rect 8356 24572 8362 24573
rect 8250 24558 8362 24572
rect 8250 24544 8264 24558
rect 8356 24556 8362 24558
rect 8379 24556 8385 24573
rect 8356 24553 8385 24556
rect 11305 24573 11326 24576
rect 11305 24556 11311 24573
rect 11305 24553 11326 24556
rect 11323 24552 11326 24553
rect 11352 24552 11355 24578
rect 13310 24572 13324 24587
rect 13807 24586 13810 24592
rect 13836 24586 13839 24612
rect 13946 24607 13975 24610
rect 13946 24590 13952 24607
rect 13969 24606 13975 24607
rect 13991 24606 13994 24612
rect 13969 24592 13994 24606
rect 13969 24590 13975 24592
rect 13946 24587 13975 24590
rect 13991 24586 13994 24592
rect 14020 24586 14023 24612
rect 14038 24607 14067 24610
rect 14038 24590 14044 24607
rect 14061 24606 14067 24607
rect 14497 24606 14500 24612
rect 14061 24592 14500 24606
rect 14061 24590 14067 24592
rect 14038 24587 14067 24590
rect 14497 24586 14500 24592
rect 14526 24606 14529 24612
rect 14819 24606 14822 24612
rect 14526 24592 14822 24606
rect 14526 24586 14529 24592
rect 14819 24586 14822 24592
rect 14848 24586 14851 24612
rect 14865 24586 14868 24612
rect 14894 24586 14897 24612
rect 16705 24586 16708 24612
rect 16734 24586 16737 24612
rect 16944 24610 16958 24626
rect 17257 24620 17260 24626
rect 17286 24620 17289 24646
rect 18591 24620 18594 24646
rect 18620 24620 18623 24646
rect 19419 24620 19422 24646
rect 19448 24640 19451 24646
rect 21903 24640 21906 24646
rect 19448 24626 19626 24640
rect 19448 24620 19451 24626
rect 16936 24607 16965 24610
rect 16936 24590 16942 24607
rect 16959 24590 16965 24607
rect 16936 24587 16965 24590
rect 17073 24586 17076 24612
rect 17102 24586 17105 24612
rect 17212 24607 17241 24610
rect 17212 24590 17218 24607
rect 17235 24606 17241 24607
rect 17901 24606 17904 24612
rect 17235 24592 17904 24606
rect 17235 24590 17241 24592
rect 17212 24587 17241 24590
rect 17901 24586 17904 24592
rect 17930 24586 17933 24612
rect 18545 24586 18548 24612
rect 18574 24586 18577 24612
rect 19557 24586 19560 24612
rect 19586 24586 19589 24612
rect 19612 24606 19626 24626
rect 20693 24626 21906 24640
rect 19757 24607 19786 24610
rect 19757 24606 19763 24607
rect 19612 24592 19763 24606
rect 19757 24590 19763 24592
rect 19780 24606 19786 24607
rect 20247 24606 20250 24612
rect 19780 24592 20250 24606
rect 19780 24590 19786 24592
rect 19757 24587 19786 24590
rect 20247 24586 20250 24592
rect 20276 24606 20279 24612
rect 20693 24606 20707 24626
rect 21903 24620 21906 24626
rect 21932 24640 21935 24646
rect 21932 24626 22018 24640
rect 21932 24620 21935 24626
rect 20276 24592 20707 24606
rect 20276 24586 20279 24592
rect 21673 24586 21676 24612
rect 21702 24606 21705 24612
rect 21950 24607 21979 24610
rect 21950 24606 21956 24607
rect 21702 24592 21956 24606
rect 21702 24586 21705 24592
rect 21950 24590 21956 24592
rect 21973 24590 21979 24607
rect 22004 24606 22018 24626
rect 22004 24592 22202 24606
rect 21950 24587 21979 24590
rect 14874 24572 14888 24586
rect 13310 24558 14888 24572
rect 15647 24552 15650 24578
rect 15676 24572 15679 24578
rect 15740 24573 15769 24576
rect 15740 24572 15746 24573
rect 15676 24558 15746 24572
rect 15676 24552 15679 24558
rect 15740 24556 15746 24558
rect 15763 24572 15769 24573
rect 15763 24558 15877 24572
rect 15763 24556 15769 24558
rect 15740 24553 15769 24556
rect 8057 24538 8060 24544
rect 7836 24524 8060 24538
rect 8057 24518 8060 24524
rect 8086 24518 8089 24544
rect 8241 24518 8244 24544
rect 8270 24518 8273 24544
rect 9231 24539 9260 24542
rect 9231 24522 9237 24539
rect 9254 24538 9260 24539
rect 9299 24538 9302 24544
rect 9254 24524 9302 24538
rect 9254 24522 9260 24524
rect 9231 24519 9260 24522
rect 9299 24518 9302 24524
rect 9328 24518 9331 24544
rect 10679 24518 10682 24544
rect 10708 24538 10711 24544
rect 12151 24542 12154 24544
rect 10726 24539 10755 24542
rect 10726 24538 10732 24539
rect 10708 24524 10732 24538
rect 10708 24518 10711 24524
rect 10726 24522 10732 24524
rect 10749 24522 10755 24539
rect 10726 24519 10755 24522
rect 12129 24539 12154 24542
rect 12129 24522 12135 24539
rect 12152 24522 12154 24539
rect 12129 24519 12154 24522
rect 12151 24518 12154 24519
rect 12180 24518 12183 24544
rect 12795 24518 12798 24544
rect 12824 24538 12827 24544
rect 13072 24539 13101 24542
rect 13072 24538 13078 24539
rect 12824 24524 13078 24538
rect 12824 24518 12827 24524
rect 13072 24522 13078 24524
rect 13095 24522 13101 24539
rect 13072 24519 13101 24522
rect 13669 24518 13672 24544
rect 13698 24518 13701 24544
rect 14866 24539 14895 24542
rect 14866 24522 14872 24539
rect 14889 24538 14895 24539
rect 15049 24538 15052 24544
rect 14889 24524 15052 24538
rect 14889 24522 14895 24524
rect 14866 24519 14895 24522
rect 15049 24518 15052 24524
rect 15078 24518 15081 24544
rect 15863 24538 15877 24558
rect 19603 24552 19606 24578
rect 19632 24572 19635 24578
rect 19718 24573 19747 24576
rect 19718 24572 19724 24573
rect 19632 24558 19724 24572
rect 19632 24552 19635 24558
rect 19718 24556 19724 24558
rect 19741 24556 19747 24573
rect 19718 24553 19747 24556
rect 21995 24552 21998 24578
rect 22024 24572 22027 24578
rect 22188 24576 22202 24592
rect 23927 24586 23930 24612
rect 23956 24606 23959 24612
rect 23974 24607 24003 24610
rect 23974 24606 23980 24607
rect 23956 24592 23980 24606
rect 23956 24586 23959 24592
rect 23974 24590 23980 24592
rect 23997 24590 24003 24607
rect 23974 24587 24003 24590
rect 22110 24573 22139 24576
rect 22110 24572 22116 24573
rect 22024 24558 22116 24572
rect 22024 24552 22027 24558
rect 22110 24556 22116 24558
rect 22133 24556 22139 24573
rect 22110 24553 22139 24556
rect 22161 24573 22202 24576
rect 22161 24556 22167 24573
rect 22184 24558 22202 24573
rect 22184 24556 22190 24558
rect 22161 24553 22190 24556
rect 24065 24552 24068 24578
rect 24094 24552 24097 24578
rect 16614 24539 16643 24542
rect 16614 24538 16620 24539
rect 15863 24524 16620 24538
rect 16614 24522 16620 24524
rect 16637 24522 16643 24539
rect 16614 24519 16643 24522
rect 20385 24518 20388 24544
rect 20414 24538 20417 24544
rect 20593 24539 20622 24542
rect 20593 24538 20599 24539
rect 20414 24524 20599 24538
rect 20414 24518 20417 24524
rect 20593 24522 20599 24524
rect 20616 24522 20622 24539
rect 20593 24519 20622 24522
rect 3036 24456 29992 24504
rect 7735 24416 7738 24442
rect 7764 24436 7767 24442
rect 7943 24437 7972 24440
rect 7943 24436 7949 24437
rect 7764 24422 7949 24436
rect 7764 24416 7767 24422
rect 7943 24420 7949 24422
rect 7966 24420 7972 24437
rect 7943 24417 7972 24420
rect 8011 24416 8014 24442
rect 8040 24436 8043 24442
rect 10725 24436 10728 24442
rect 8040 24422 10728 24436
rect 8040 24416 8043 24422
rect 10725 24416 10728 24422
rect 10754 24436 10757 24442
rect 12105 24436 12108 24442
rect 10754 24422 12108 24436
rect 10754 24416 10757 24422
rect 12105 24416 12108 24422
rect 12134 24416 12137 24442
rect 13991 24416 13994 24442
rect 14020 24436 14023 24442
rect 14175 24436 14178 24442
rect 14020 24422 14178 24436
rect 14020 24416 14023 24422
rect 14175 24416 14178 24422
rect 14204 24436 14207 24442
rect 16153 24436 16156 24442
rect 14204 24422 16156 24436
rect 14204 24416 14207 24422
rect 16153 24416 16156 24422
rect 16182 24416 16185 24442
rect 17763 24416 17766 24442
rect 17792 24416 17795 24442
rect 21075 24436 21078 24442
rect 20348 24422 20868 24436
rect 8057 24382 8060 24408
rect 8086 24402 8089 24408
rect 8086 24388 9276 24402
rect 8086 24382 8089 24388
rect 9262 24374 9276 24388
rect 9299 24382 9302 24408
rect 9328 24382 9331 24408
rect 12427 24402 12430 24408
rect 12283 24388 12430 24402
rect 3273 24348 3276 24374
rect 3302 24368 3305 24374
rect 3503 24368 3506 24374
rect 3302 24354 3506 24368
rect 3302 24348 3305 24354
rect 3503 24348 3506 24354
rect 3532 24368 3535 24374
rect 3613 24369 3642 24372
rect 3613 24368 3619 24369
rect 3532 24354 3619 24368
rect 3532 24348 3535 24354
rect 3613 24352 3619 24354
rect 3636 24352 3642 24369
rect 3613 24349 3642 24352
rect 3657 24369 3686 24372
rect 3657 24352 3663 24369
rect 3680 24368 3686 24369
rect 5849 24368 5852 24374
rect 3680 24354 5852 24368
rect 3680 24352 3686 24354
rect 3657 24349 3686 24352
rect 5849 24348 5852 24354
rect 5878 24348 5881 24374
rect 7045 24348 7048 24374
rect 7074 24372 7077 24374
rect 7074 24369 7092 24372
rect 7086 24352 7092 24369
rect 7074 24349 7092 24352
rect 7107 24369 7136 24372
rect 7107 24352 7113 24369
rect 7130 24368 7136 24369
rect 7551 24368 7554 24374
rect 7130 24354 7554 24368
rect 7130 24352 7136 24354
rect 7107 24349 7136 24352
rect 7074 24348 7077 24349
rect 7551 24348 7554 24354
rect 7580 24348 7583 24374
rect 9161 24348 9164 24374
rect 9190 24348 9193 24374
rect 9253 24348 9256 24374
rect 9282 24348 9285 24374
rect 9345 24348 9348 24374
rect 9374 24372 9377 24374
rect 9374 24368 9378 24372
rect 9374 24354 9396 24368
rect 9374 24349 9378 24354
rect 9374 24348 9377 24349
rect 10541 24348 10544 24374
rect 10570 24368 10573 24374
rect 12013 24368 12016 24374
rect 10570 24354 12016 24368
rect 10570 24348 10573 24354
rect 12013 24348 12016 24354
rect 12042 24348 12045 24374
rect 12059 24348 12062 24374
rect 12088 24372 12091 24374
rect 12088 24369 12100 24372
rect 12094 24352 12100 24369
rect 12088 24349 12100 24352
rect 12088 24348 12091 24349
rect 12151 24348 12154 24374
rect 12180 24372 12183 24374
rect 12180 24369 12194 24372
rect 12188 24352 12194 24369
rect 12283 24367 12297 24388
rect 12427 24382 12430 24388
rect 12456 24382 12459 24408
rect 14911 24382 14914 24408
rect 14940 24402 14943 24408
rect 16015 24402 16018 24408
rect 14940 24388 16018 24402
rect 14940 24382 14943 24388
rect 16015 24382 16018 24388
rect 16044 24402 16047 24408
rect 16044 24388 16360 24402
rect 16044 24382 16047 24388
rect 12335 24372 12338 24374
rect 12326 24369 12338 24372
rect 12180 24349 12194 24352
rect 12227 24364 12256 24367
rect 12180 24348 12183 24349
rect 12227 24347 12233 24364
rect 12250 24347 12256 24364
rect 12227 24344 12256 24347
rect 12275 24364 12304 24367
rect 12275 24347 12281 24364
rect 12298 24347 12304 24364
rect 12326 24352 12332 24369
rect 12364 24368 12367 24374
rect 15141 24368 15144 24374
rect 12364 24354 15144 24368
rect 12326 24349 12338 24352
rect 12335 24348 12338 24349
rect 12364 24348 12367 24354
rect 15141 24348 15144 24354
rect 15170 24348 15173 24374
rect 16062 24369 16091 24372
rect 16062 24352 16068 24369
rect 16085 24352 16091 24369
rect 16062 24349 16091 24352
rect 12275 24344 12304 24347
rect 3411 24314 3414 24340
rect 3440 24334 3443 24340
rect 3458 24335 3487 24338
rect 3458 24334 3464 24335
rect 3440 24320 3464 24334
rect 3440 24314 3443 24320
rect 3458 24318 3464 24320
rect 3481 24318 3487 24335
rect 3458 24315 3487 24318
rect 6907 24314 6910 24340
rect 6936 24314 6939 24340
rect 9300 24335 9329 24338
rect 9300 24318 9306 24335
rect 9323 24334 9329 24335
rect 9437 24334 9440 24340
rect 9323 24320 9440 24334
rect 9323 24318 9329 24320
rect 9300 24315 9329 24318
rect 9437 24314 9440 24320
rect 9466 24314 9469 24340
rect 12235 24300 12249 24344
rect 13807 24314 13810 24340
rect 13836 24334 13839 24340
rect 13991 24334 13994 24340
rect 13836 24320 13994 24334
rect 13836 24314 13839 24320
rect 13991 24314 13994 24320
rect 14020 24334 14023 24340
rect 14451 24334 14454 24340
rect 14020 24320 14454 24334
rect 14020 24314 14023 24320
rect 14451 24314 14454 24320
rect 14480 24334 14483 24340
rect 16070 24334 16084 24349
rect 16153 24348 16156 24374
rect 16182 24348 16185 24374
rect 16346 24372 16360 24388
rect 16338 24369 16367 24372
rect 16338 24352 16344 24369
rect 16361 24352 16367 24369
rect 17580 24369 17609 24372
rect 17580 24368 17586 24369
rect 16338 24349 16367 24352
rect 16392 24354 17586 24368
rect 16392 24334 16406 24354
rect 17580 24352 17586 24354
rect 17603 24368 17609 24369
rect 17717 24368 17720 24374
rect 17603 24354 17720 24368
rect 17603 24352 17609 24354
rect 17580 24349 17609 24352
rect 17717 24348 17720 24354
rect 17746 24348 17749 24374
rect 19603 24348 19606 24374
rect 19632 24368 19635 24374
rect 20348 24372 20362 24422
rect 20340 24369 20369 24372
rect 20340 24368 20346 24369
rect 19632 24354 20346 24368
rect 19632 24348 19635 24354
rect 20340 24352 20346 24354
rect 20363 24352 20369 24369
rect 20754 24369 20783 24372
rect 20754 24368 20760 24369
rect 20340 24349 20369 24352
rect 20532 24354 20760 24368
rect 14480 24320 16406 24334
rect 14480 24314 14483 24320
rect 17533 24314 17536 24340
rect 17562 24314 17565 24340
rect 20385 24314 20388 24340
rect 20414 24314 20417 24340
rect 20532 24338 20546 24354
rect 20754 24352 20760 24354
rect 20777 24352 20783 24369
rect 20754 24349 20783 24352
rect 20524 24335 20553 24338
rect 20524 24318 20530 24335
rect 20547 24318 20553 24335
rect 20854 24334 20868 24422
rect 20900 24422 21078 24436
rect 20900 24372 20914 24422
rect 21075 24416 21078 24422
rect 21104 24416 21107 24442
rect 23422 24437 23451 24440
rect 23422 24420 23428 24437
rect 23445 24436 23451 24437
rect 23559 24436 23562 24442
rect 23445 24422 23562 24436
rect 23445 24420 23451 24422
rect 23422 24417 23451 24420
rect 23559 24416 23562 24422
rect 23588 24416 23591 24442
rect 22823 24402 22826 24408
rect 20946 24388 22826 24402
rect 20892 24369 20921 24372
rect 20892 24352 20898 24369
rect 20915 24352 20921 24369
rect 20892 24349 20921 24352
rect 20946 24334 20960 24388
rect 22823 24382 22826 24388
rect 22852 24382 22855 24408
rect 22878 24388 23444 24402
rect 20983 24348 20986 24374
rect 21012 24348 21015 24374
rect 21122 24369 21151 24372
rect 21122 24352 21128 24369
rect 21145 24352 21151 24369
rect 21122 24349 21151 24352
rect 20854 24320 20960 24334
rect 20524 24315 20553 24318
rect 12381 24300 12384 24306
rect 12235 24286 12384 24300
rect 12381 24280 12384 24286
rect 12410 24280 12413 24306
rect 16337 24280 16340 24306
rect 16366 24280 16369 24306
rect 4493 24267 4522 24270
rect 4493 24250 4499 24267
rect 4516 24266 4522 24267
rect 5021 24266 5024 24272
rect 4516 24252 5024 24266
rect 4516 24250 4522 24252
rect 4493 24247 4522 24250
rect 5021 24246 5024 24252
rect 5050 24246 5053 24272
rect 6493 24246 6496 24272
rect 6522 24266 6525 24272
rect 9345 24266 9348 24272
rect 6522 24252 9348 24266
rect 6522 24246 6525 24252
rect 9345 24246 9348 24252
rect 9374 24266 9377 24272
rect 9621 24266 9624 24272
rect 9374 24252 9624 24266
rect 9374 24246 9377 24252
rect 9621 24246 9624 24252
rect 9650 24246 9653 24272
rect 12014 24267 12043 24270
rect 12014 24250 12020 24267
rect 12037 24266 12043 24267
rect 12151 24266 12154 24272
rect 12037 24252 12154 24266
rect 12037 24250 12043 24252
rect 12014 24247 12043 24250
rect 12151 24246 12154 24252
rect 12180 24246 12183 24272
rect 21130 24266 21144 24349
rect 22087 24348 22090 24374
rect 22116 24368 22119 24374
rect 22878 24368 22892 24388
rect 22116 24354 22892 24368
rect 22116 24348 22119 24354
rect 22961 24348 22964 24374
rect 22990 24368 22993 24374
rect 23237 24368 23240 24374
rect 22990 24354 23240 24368
rect 22990 24348 22993 24354
rect 23237 24348 23240 24354
rect 23266 24348 23269 24374
rect 23375 24348 23378 24374
rect 23404 24348 23407 24374
rect 23430 24368 23444 24388
rect 23467 24382 23470 24408
rect 23496 24406 23499 24408
rect 23496 24403 23507 24406
rect 23501 24386 23507 24403
rect 24111 24402 24114 24408
rect 23496 24383 23507 24386
rect 23614 24388 24114 24402
rect 23496 24382 23499 24383
rect 23614 24368 23628 24388
rect 24111 24382 24114 24388
rect 24140 24402 24143 24408
rect 24296 24403 24325 24406
rect 24296 24402 24302 24403
rect 24140 24388 24302 24402
rect 24140 24382 24143 24388
rect 24296 24386 24302 24388
rect 24319 24386 24325 24403
rect 24296 24383 24325 24386
rect 23430 24354 23628 24368
rect 23743 24348 23746 24374
rect 23772 24368 23775 24374
rect 23928 24369 23957 24372
rect 23928 24368 23934 24369
rect 23772 24354 23934 24368
rect 23772 24348 23775 24354
rect 23928 24352 23934 24354
rect 23951 24352 23957 24369
rect 23928 24349 23957 24352
rect 24020 24369 24049 24372
rect 24020 24352 24026 24369
rect 24043 24352 24049 24369
rect 24020 24349 24049 24352
rect 21167 24314 21170 24340
rect 21196 24314 21199 24340
rect 22915 24314 22918 24340
rect 22944 24314 22947 24340
rect 23560 24335 23589 24338
rect 23560 24334 23566 24335
rect 23154 24320 23566 24334
rect 23154 24304 23168 24320
rect 23560 24318 23566 24320
rect 23583 24318 23589 24335
rect 24028 24334 24042 24349
rect 24065 24348 24068 24374
rect 24094 24348 24097 24374
rect 24111 24334 24114 24340
rect 24028 24320 24114 24334
rect 23560 24315 23589 24318
rect 24111 24314 24114 24320
rect 24140 24314 24143 24340
rect 23146 24301 23175 24304
rect 23146 24284 23152 24301
rect 23169 24284 23175 24301
rect 23146 24281 23175 24284
rect 23283 24280 23286 24306
rect 23312 24300 23315 24306
rect 24342 24301 24371 24304
rect 24342 24300 24348 24301
rect 23312 24286 24348 24300
rect 23312 24280 23315 24286
rect 24342 24284 24348 24286
rect 24365 24300 24371 24301
rect 24617 24300 24620 24306
rect 24365 24286 24620 24300
rect 24365 24284 24371 24286
rect 24342 24281 24371 24284
rect 24617 24280 24620 24286
rect 24646 24280 24649 24306
rect 23422 24267 23451 24270
rect 23422 24266 23428 24267
rect 21130 24252 23428 24266
rect 23422 24250 23428 24252
rect 23445 24250 23451 24267
rect 23422 24247 23451 24250
rect 23927 24246 23930 24272
rect 23956 24246 23959 24272
rect 3036 24184 29992 24232
rect 3411 24164 3414 24170
rect 3144 24150 3414 24164
rect 3144 24100 3158 24150
rect 3411 24144 3414 24150
rect 3440 24144 3443 24170
rect 8195 24164 8198 24170
rect 8066 24150 8198 24164
rect 5022 24131 5051 24134
rect 5022 24114 5028 24131
rect 5045 24130 5051 24131
rect 5067 24130 5070 24136
rect 5045 24116 5070 24130
rect 5045 24114 5051 24116
rect 5022 24111 5051 24114
rect 5067 24110 5070 24116
rect 5096 24110 5099 24136
rect 5527 24110 5530 24136
rect 5556 24130 5559 24136
rect 5665 24130 5668 24136
rect 5556 24116 5668 24130
rect 5556 24110 5559 24116
rect 5665 24110 5668 24116
rect 5694 24130 5697 24136
rect 7045 24130 7048 24136
rect 5694 24116 7048 24130
rect 5694 24110 5697 24116
rect 7045 24110 7048 24116
rect 7074 24110 7077 24136
rect 3136 24097 3165 24100
rect 3136 24080 3142 24097
rect 3159 24080 3165 24097
rect 3136 24077 3165 24080
rect 6907 24076 6910 24102
rect 6936 24096 6939 24102
rect 8066 24100 8080 24150
rect 8195 24144 8198 24150
rect 8224 24164 8227 24170
rect 9093 24165 9122 24168
rect 8224 24150 9000 24164
rect 8224 24144 8227 24150
rect 8986 24130 9000 24150
rect 9093 24148 9099 24165
rect 9116 24164 9122 24165
rect 9161 24164 9164 24170
rect 9116 24150 9164 24164
rect 9116 24148 9122 24150
rect 9093 24145 9122 24148
rect 9161 24144 9164 24150
rect 9190 24144 9193 24170
rect 9207 24144 9210 24170
rect 9236 24164 9239 24170
rect 13209 24164 13212 24170
rect 9236 24150 13212 24164
rect 9236 24144 9239 24150
rect 13209 24144 13212 24150
rect 13238 24164 13241 24170
rect 13669 24164 13672 24170
rect 13238 24150 13672 24164
rect 13238 24144 13241 24150
rect 13669 24144 13672 24150
rect 13698 24144 13701 24170
rect 22755 24165 22784 24168
rect 22755 24148 22761 24165
rect 22778 24164 22784 24165
rect 22915 24164 22918 24170
rect 22778 24150 22918 24164
rect 22778 24148 22784 24150
rect 22755 24145 22784 24148
rect 22915 24144 22918 24150
rect 22944 24144 22947 24170
rect 9023 24130 9026 24136
rect 8986 24116 9026 24130
rect 9023 24110 9026 24116
rect 9052 24110 9055 24136
rect 15863 24116 17234 24130
rect 8058 24097 8087 24100
rect 8058 24096 8064 24097
rect 6936 24082 8064 24096
rect 6936 24076 6939 24082
rect 8058 24080 8064 24082
rect 8081 24080 8087 24097
rect 8058 24077 8087 24080
rect 12336 24097 12365 24100
rect 12336 24080 12342 24097
rect 12359 24096 12365 24097
rect 15863 24096 15877 24116
rect 12359 24082 15877 24096
rect 12359 24080 12365 24082
rect 12336 24077 12365 24080
rect 16291 24076 16294 24102
rect 16320 24096 16323 24102
rect 17074 24097 17103 24100
rect 17074 24096 17080 24097
rect 16320 24082 17080 24096
rect 16320 24076 16323 24082
rect 17074 24080 17080 24082
rect 17097 24096 17103 24097
rect 17119 24096 17122 24102
rect 17097 24082 17122 24096
rect 17097 24080 17103 24082
rect 17074 24077 17103 24080
rect 17119 24076 17122 24082
rect 17148 24076 17151 24102
rect 17220 24096 17234 24116
rect 18453 24110 18456 24136
rect 18482 24110 18485 24136
rect 20662 24131 20691 24134
rect 20662 24114 20668 24131
rect 20685 24130 20691 24131
rect 20983 24130 20986 24136
rect 20685 24116 20986 24130
rect 20685 24114 20691 24116
rect 20662 24111 20691 24114
rect 20983 24110 20986 24116
rect 21012 24110 21015 24136
rect 24433 24110 24436 24136
rect 24462 24130 24465 24136
rect 24480 24131 24509 24134
rect 24480 24130 24486 24131
rect 24462 24116 24486 24130
rect 24462 24110 24465 24116
rect 24480 24114 24486 24116
rect 24503 24114 24509 24131
rect 24480 24111 24509 24114
rect 18637 24096 18640 24102
rect 17220 24082 18640 24096
rect 18637 24076 18640 24082
rect 18666 24076 18669 24102
rect 20431 24076 20434 24102
rect 20460 24076 20463 24102
rect 21673 24076 21676 24102
rect 21702 24096 21705 24102
rect 21720 24097 21749 24100
rect 21720 24096 21726 24097
rect 21702 24082 21726 24096
rect 21702 24076 21705 24082
rect 21720 24080 21726 24082
rect 21743 24080 21749 24097
rect 21720 24077 21749 24080
rect 24249 24076 24252 24102
rect 24278 24076 24281 24102
rect 3297 24063 3326 24066
rect 3297 24046 3303 24063
rect 3320 24062 3326 24063
rect 3457 24062 3460 24068
rect 3320 24048 3460 24062
rect 3320 24046 3326 24048
rect 3297 24043 3326 24046
rect 3457 24042 3460 24048
rect 3486 24042 3489 24068
rect 4929 24042 4932 24068
rect 4958 24062 4961 24068
rect 5114 24063 5143 24066
rect 5114 24062 5120 24063
rect 4958 24048 5120 24062
rect 4958 24042 4961 24048
rect 5114 24046 5120 24048
rect 5137 24046 5143 24063
rect 5114 24043 5143 24046
rect 8219 24063 8248 24066
rect 8219 24046 8225 24063
rect 8242 24062 8248 24063
rect 8333 24062 8336 24068
rect 8242 24048 8336 24062
rect 8242 24046 8248 24048
rect 8219 24043 8248 24046
rect 8333 24042 8336 24048
rect 8362 24062 8365 24068
rect 9161 24062 9164 24068
rect 8362 24048 9164 24062
rect 8362 24042 8365 24048
rect 9161 24042 9164 24048
rect 9190 24042 9193 24068
rect 12151 24042 12154 24068
rect 12180 24042 12183 24068
rect 12289 24042 12292 24068
rect 12318 24042 12321 24068
rect 12382 24063 12411 24066
rect 12382 24046 12388 24063
rect 12405 24062 12411 24063
rect 12657 24062 12660 24068
rect 12405 24048 12660 24062
rect 12405 24046 12411 24048
rect 12382 24043 12411 24046
rect 12657 24042 12660 24048
rect 12686 24042 12689 24068
rect 13991 24042 13994 24068
rect 14020 24042 14023 24068
rect 14175 24042 14178 24068
rect 14204 24042 14207 24068
rect 14268 24063 14297 24066
rect 14268 24046 14274 24063
rect 14291 24062 14297 24063
rect 14497 24062 14500 24068
rect 14291 24048 14500 24062
rect 14291 24046 14297 24048
rect 14268 24043 14297 24046
rect 14497 24042 14500 24048
rect 14526 24062 14529 24068
rect 14865 24062 14868 24068
rect 14526 24048 14868 24062
rect 14526 24042 14529 24048
rect 14865 24042 14868 24048
rect 14894 24042 14897 24068
rect 16337 24042 16340 24068
rect 16366 24042 16369 24068
rect 16705 24042 16708 24068
rect 16734 24062 16737 24068
rect 16844 24063 16873 24066
rect 16844 24062 16850 24063
rect 16734 24048 16850 24062
rect 16734 24042 16737 24048
rect 16844 24046 16850 24048
rect 16867 24046 16873 24063
rect 16844 24043 16873 24046
rect 17028 24063 17057 24066
rect 17028 24046 17034 24063
rect 17051 24062 17057 24063
rect 17901 24062 17904 24068
rect 17051 24048 17904 24062
rect 17051 24046 17057 24048
rect 17028 24043 17057 24046
rect 17901 24042 17904 24048
rect 17930 24042 17933 24068
rect 18085 24042 18088 24068
rect 18114 24062 18117 24068
rect 18591 24062 18594 24068
rect 18114 24048 18594 24062
rect 18114 24042 18117 24048
rect 18591 24042 18594 24048
rect 18620 24042 18623 24068
rect 20017 24042 20020 24068
rect 20046 24062 20049 24068
rect 20478 24063 20507 24066
rect 20478 24062 20484 24063
rect 20046 24048 20484 24062
rect 20046 24042 20049 24048
rect 20478 24046 20484 24048
rect 20501 24046 20507 24063
rect 20478 24043 20507 24046
rect 21397 24042 21400 24068
rect 21426 24062 21429 24068
rect 21881 24063 21910 24066
rect 21881 24062 21887 24063
rect 21426 24048 21887 24062
rect 21426 24042 21429 24048
rect 21881 24046 21887 24048
rect 21904 24062 21910 24063
rect 23237 24062 23240 24068
rect 21904 24048 23240 24062
rect 21904 24046 21910 24048
rect 21881 24043 21910 24046
rect 23237 24042 23240 24048
rect 23266 24042 23269 24068
rect 24111 24042 24114 24068
rect 24140 24042 24143 24068
rect 24158 24063 24187 24066
rect 24158 24046 24164 24063
rect 24181 24062 24187 24063
rect 24181 24048 24594 24062
rect 24181 24046 24187 24048
rect 24158 24043 24187 24046
rect 3181 24008 3184 24034
rect 3210 24028 3213 24034
rect 3365 24032 3368 24034
rect 3347 24029 3368 24032
rect 3347 24028 3353 24029
rect 3210 24014 3353 24028
rect 3210 24008 3213 24014
rect 3347 24012 3353 24014
rect 3347 24009 3368 24012
rect 3365 24008 3368 24009
rect 3394 24008 3397 24034
rect 4976 24029 5005 24032
rect 4976 24012 4982 24029
rect 4999 24012 5005 24029
rect 4976 24009 5005 24012
rect 5068 24029 5097 24032
rect 5068 24012 5074 24029
rect 5091 24028 5097 24029
rect 6953 24028 6956 24034
rect 5091 24014 6956 24028
rect 5091 24012 5097 24014
rect 5068 24009 5097 24012
rect 4171 23995 4200 23998
rect 4171 23978 4177 23995
rect 4194 23994 4200 23995
rect 4745 23994 4748 24000
rect 4194 23980 4748 23994
rect 4194 23978 4200 23980
rect 4171 23975 4200 23978
rect 4745 23974 4748 23980
rect 4774 23974 4777 24000
rect 4984 23994 4998 24009
rect 6953 24008 6956 24014
rect 6982 24008 6985 24034
rect 7551 24008 7554 24034
rect 7580 24028 7583 24034
rect 8265 24029 8294 24032
rect 8265 24028 8271 24029
rect 7580 24014 8271 24028
rect 7580 24008 7583 24014
rect 8265 24012 8271 24014
rect 8288 24012 8294 24029
rect 8265 24009 8294 24012
rect 18454 24029 18483 24032
rect 18454 24012 18460 24029
rect 18477 24028 18483 24029
rect 18499 24028 18502 24034
rect 18477 24014 18502 24028
rect 18477 24012 18483 24014
rect 18454 24009 18483 24012
rect 18499 24008 18502 24014
rect 18528 24008 18531 24034
rect 21949 24032 21952 24034
rect 21931 24029 21952 24032
rect 21931 24012 21937 24029
rect 21931 24009 21952 24012
rect 21949 24008 21952 24009
rect 21978 24008 21981 24034
rect 24250 24029 24279 24032
rect 24250 24012 24256 24029
rect 24273 24028 24279 24029
rect 24480 24029 24509 24032
rect 24480 24028 24486 24029
rect 24273 24014 24486 24028
rect 24273 24012 24279 24014
rect 24250 24009 24279 24012
rect 24480 24012 24486 24014
rect 24503 24012 24509 24029
rect 24580 24028 24594 24048
rect 24617 24042 24620 24068
rect 24646 24042 24649 24068
rect 24801 24028 24804 24034
rect 24580 24014 24804 24028
rect 24480 24009 24509 24012
rect 24801 24008 24804 24014
rect 24830 24008 24833 24034
rect 5573 23994 5576 24000
rect 4984 23980 5576 23994
rect 5573 23974 5576 23980
rect 5602 23974 5605 24000
rect 13899 23974 13902 24000
rect 13928 23974 13931 24000
rect 16383 23974 16386 24000
rect 16412 23974 16415 24000
rect 16982 23995 17011 23998
rect 16982 23978 16988 23995
rect 17005 23994 17011 23995
rect 17027 23994 17030 24000
rect 17005 23980 17030 23994
rect 17005 23978 17011 23980
rect 16982 23975 17011 23978
rect 17027 23974 17030 23980
rect 17056 23974 17059 24000
rect 17993 23974 17996 24000
rect 18022 23994 18025 24000
rect 18546 23995 18575 23998
rect 18546 23994 18552 23995
rect 18022 23980 18552 23994
rect 18022 23974 18025 23980
rect 18546 23978 18552 23980
rect 18569 23994 18575 23995
rect 18591 23994 18594 24000
rect 18569 23980 18594 23994
rect 18569 23978 18575 23980
rect 18546 23975 18575 23978
rect 18591 23974 18594 23980
rect 18620 23974 18623 24000
rect 23605 23974 23608 24000
rect 23634 23994 23637 24000
rect 24111 23994 24114 24000
rect 23634 23980 24114 23994
rect 23634 23974 23637 23980
rect 24111 23974 24114 23980
rect 24140 23994 24143 24000
rect 24572 23995 24601 23998
rect 24572 23994 24578 23995
rect 24140 23980 24578 23994
rect 24140 23974 24143 23980
rect 24572 23978 24578 23980
rect 24595 23978 24601 23995
rect 24572 23975 24601 23978
rect 3036 23912 29992 23960
rect 4837 23892 4840 23898
rect 4823 23872 4840 23892
rect 4866 23872 4869 23898
rect 4929 23872 4932 23898
rect 4958 23892 4961 23898
rect 4976 23893 5005 23896
rect 4976 23892 4982 23893
rect 4958 23878 4982 23892
rect 4958 23872 4961 23878
rect 4976 23876 4982 23878
rect 4999 23876 5005 23893
rect 4976 23873 5005 23876
rect 5021 23872 5024 23898
rect 5050 23872 5053 23898
rect 17901 23872 17904 23898
rect 17930 23892 17933 23898
rect 19006 23893 19035 23896
rect 19006 23892 19012 23893
rect 17930 23878 19012 23892
rect 17930 23872 17933 23878
rect 19006 23876 19012 23878
rect 19029 23876 19035 23893
rect 19006 23873 19035 23876
rect 21398 23893 21427 23896
rect 21398 23876 21404 23893
rect 21421 23892 21427 23893
rect 21581 23892 21584 23898
rect 21421 23878 21584 23892
rect 21421 23876 21427 23878
rect 21398 23873 21427 23876
rect 21581 23872 21584 23878
rect 21610 23872 21613 23898
rect 23743 23872 23746 23898
rect 23772 23872 23775 23898
rect 24249 23892 24252 23898
rect 23890 23878 24252 23892
rect 3457 23838 3460 23864
rect 3486 23858 3489 23864
rect 3687 23862 3690 23864
rect 3618 23859 3647 23862
rect 3618 23858 3624 23859
rect 3486 23844 3624 23858
rect 3486 23838 3489 23844
rect 3618 23842 3624 23844
rect 3641 23842 3647 23859
rect 3618 23839 3647 23842
rect 3669 23859 3690 23862
rect 3669 23842 3675 23859
rect 3669 23839 3690 23842
rect 3687 23838 3690 23839
rect 3716 23838 3719 23864
rect 4823 23858 4837 23872
rect 4800 23844 4837 23858
rect 4745 23804 4748 23830
rect 4774 23804 4777 23830
rect 4800 23828 4814 23844
rect 5030 23828 5044 23872
rect 6355 23838 6358 23864
rect 6384 23838 6387 23864
rect 6953 23838 6956 23864
rect 6982 23858 6985 23864
rect 7107 23859 7136 23862
rect 7107 23858 7113 23859
rect 6982 23844 7113 23858
rect 6982 23838 6985 23844
rect 7107 23842 7113 23844
rect 7130 23842 7136 23859
rect 13117 23858 13120 23864
rect 7107 23839 7136 23842
rect 7928 23844 9244 23858
rect 4800 23825 4842 23828
rect 4800 23810 4819 23825
rect 4813 23808 4819 23810
rect 4836 23808 4842 23825
rect 4904 23825 4933 23828
rect 4904 23824 4910 23825
rect 4813 23805 4842 23808
rect 4872 23810 4910 23824
rect 3411 23770 3414 23796
rect 3440 23790 3443 23796
rect 3458 23791 3487 23794
rect 3458 23790 3464 23791
rect 3440 23776 3464 23790
rect 3440 23770 3443 23776
rect 3458 23774 3464 23776
rect 3481 23774 3487 23791
rect 3458 23771 3487 23774
rect 4493 23791 4522 23794
rect 4493 23774 4499 23791
rect 4516 23790 4522 23791
rect 4872 23790 4886 23810
rect 4904 23808 4910 23810
rect 4927 23808 4933 23825
rect 5007 23825 5044 23828
rect 4904 23805 4933 23808
rect 4959 23820 4988 23823
rect 4959 23803 4965 23820
rect 4982 23803 4988 23820
rect 5007 23808 5013 23825
rect 5030 23810 5044 23825
rect 5058 23825 5087 23828
rect 5030 23808 5036 23810
rect 5007 23805 5036 23808
rect 5058 23808 5064 23825
rect 5081 23824 5087 23825
rect 5081 23810 6217 23824
rect 5081 23808 5087 23810
rect 5058 23805 5087 23808
rect 4959 23800 4988 23803
rect 4516 23776 4886 23790
rect 4516 23774 4522 23776
rect 4493 23771 4522 23774
rect 4883 23736 4886 23762
rect 4912 23756 4915 23762
rect 4967 23756 4981 23800
rect 6203 23790 6217 23810
rect 6447 23804 6450 23830
rect 6476 23804 6479 23830
rect 6494 23825 6523 23828
rect 6494 23808 6500 23825
rect 6517 23824 6523 23825
rect 6815 23824 6818 23830
rect 6517 23810 6818 23824
rect 6517 23808 6523 23810
rect 6494 23805 6523 23808
rect 6815 23804 6818 23810
rect 6844 23804 6847 23830
rect 6907 23804 6910 23830
rect 6936 23804 6939 23830
rect 7045 23804 7048 23830
rect 7074 23828 7077 23830
rect 7074 23825 7097 23828
rect 7091 23824 7097 23825
rect 7321 23824 7324 23830
rect 7091 23810 7324 23824
rect 7091 23808 7097 23810
rect 7074 23805 7097 23808
rect 7074 23804 7077 23805
rect 7321 23804 7324 23810
rect 7350 23804 7353 23830
rect 7928 23824 7942 23844
rect 7836 23810 7942 23824
rect 6585 23790 6588 23796
rect 6203 23776 6588 23790
rect 6585 23770 6588 23776
rect 6614 23770 6617 23796
rect 4912 23742 4981 23756
rect 5214 23742 6930 23756
rect 4912 23736 4915 23742
rect 3641 23702 3644 23728
rect 3670 23722 3673 23728
rect 5214 23722 5228 23742
rect 3670 23708 5228 23722
rect 3670 23702 3673 23708
rect 5251 23702 5254 23728
rect 5280 23722 5283 23728
rect 6033 23722 6036 23728
rect 5280 23708 6036 23722
rect 5280 23702 5283 23708
rect 6033 23702 6036 23708
rect 6062 23702 6065 23728
rect 6355 23702 6358 23728
rect 6384 23702 6387 23728
rect 6916 23722 6930 23742
rect 7836 23722 7850 23810
rect 9023 23804 9026 23830
rect 9052 23804 9055 23830
rect 9161 23804 9164 23830
rect 9190 23828 9193 23830
rect 9230 23828 9244 23844
rect 12988 23844 13120 23858
rect 9190 23825 9208 23828
rect 9202 23808 9208 23825
rect 9190 23805 9208 23808
rect 9223 23825 9252 23828
rect 9223 23808 9229 23825
rect 9246 23824 9252 23825
rect 11323 23824 11326 23830
rect 9246 23810 11326 23824
rect 9246 23808 9252 23810
rect 9223 23805 9252 23808
rect 9190 23804 9193 23805
rect 11323 23804 11326 23810
rect 11352 23804 11355 23830
rect 12988 23828 13002 23844
rect 13117 23838 13120 23844
rect 13146 23858 13149 23864
rect 13531 23858 13534 23864
rect 13146 23844 13534 23858
rect 13146 23838 13149 23844
rect 13531 23838 13534 23844
rect 13560 23838 13563 23864
rect 12980 23825 13009 23828
rect 12980 23808 12986 23825
rect 13003 23808 13009 23825
rect 12980 23805 13009 23808
rect 13072 23825 13101 23828
rect 13072 23808 13078 23825
rect 13095 23824 13101 23825
rect 13255 23824 13258 23830
rect 13095 23810 13258 23824
rect 13095 23808 13101 23810
rect 13072 23805 13101 23808
rect 13255 23804 13258 23810
rect 13284 23824 13287 23830
rect 13284 23810 13922 23824
rect 13284 23804 13287 23810
rect 7873 23770 7876 23796
rect 7902 23790 7905 23796
rect 7943 23791 7972 23794
rect 7943 23790 7949 23791
rect 7902 23776 7949 23790
rect 7902 23770 7905 23776
rect 7943 23774 7949 23776
rect 7966 23774 7972 23791
rect 7943 23771 7972 23774
rect 13210 23791 13239 23794
rect 13210 23774 13216 23791
rect 13233 23790 13239 23791
rect 13301 23790 13304 23796
rect 13233 23776 13304 23790
rect 13233 23774 13239 23776
rect 13210 23771 13239 23774
rect 13301 23770 13304 23776
rect 13330 23770 13333 23796
rect 13908 23790 13922 23810
rect 14957 23804 14960 23830
rect 14986 23804 14989 23830
rect 15049 23804 15052 23830
rect 15078 23804 15081 23830
rect 17910 23828 17924 23872
rect 18453 23862 18456 23864
rect 18450 23858 18456 23862
rect 18433 23844 18456 23858
rect 18450 23839 18456 23844
rect 18453 23838 18456 23839
rect 18482 23838 18485 23864
rect 21306 23859 21335 23862
rect 21306 23842 21312 23859
rect 21329 23858 21335 23859
rect 21673 23858 21676 23864
rect 21329 23844 21676 23858
rect 21329 23842 21335 23844
rect 21306 23839 21335 23842
rect 21673 23838 21676 23844
rect 21702 23838 21705 23864
rect 17902 23825 17931 23828
rect 17902 23808 17908 23825
rect 17925 23808 17931 23825
rect 17902 23805 17931 23808
rect 18316 23825 18345 23828
rect 18316 23808 18322 23825
rect 18339 23824 18345 23825
rect 18361 23824 18364 23830
rect 18339 23810 18364 23824
rect 18339 23808 18345 23810
rect 18316 23805 18345 23808
rect 18361 23804 18364 23810
rect 18390 23824 18393 23830
rect 19373 23824 19376 23830
rect 18390 23810 19376 23824
rect 18390 23804 18393 23810
rect 19373 23804 19376 23810
rect 19402 23824 19405 23830
rect 19557 23824 19560 23830
rect 19402 23810 19560 23824
rect 19402 23804 19405 23810
rect 19557 23804 19560 23810
rect 19586 23804 19589 23830
rect 21443 23804 21446 23830
rect 21472 23804 21475 23830
rect 23890 23824 23904 23878
rect 24249 23872 24252 23878
rect 24278 23872 24281 23898
rect 23927 23838 23930 23864
rect 23956 23858 23959 23864
rect 24097 23859 24126 23862
rect 24097 23858 24103 23859
rect 23956 23844 24103 23858
rect 23956 23838 23959 23844
rect 24097 23842 24103 23844
rect 24120 23842 24126 23859
rect 24097 23839 24126 23842
rect 23568 23810 23904 23824
rect 23974 23825 24003 23828
rect 15058 23790 15072 23804
rect 13908 23776 15072 23790
rect 15187 23770 15190 23796
rect 15216 23770 15219 23796
rect 17947 23770 17950 23796
rect 17976 23770 17979 23796
rect 18085 23770 18088 23796
rect 18114 23770 18117 23796
rect 21305 23770 21308 23796
rect 21334 23790 21337 23796
rect 23568 23790 23582 23810
rect 21334 23776 23582 23790
rect 21334 23770 21337 23776
rect 23605 23770 23608 23796
rect 23634 23770 23637 23796
rect 23752 23794 23766 23810
rect 23974 23808 23980 23825
rect 23997 23824 24003 23825
rect 24387 23824 24390 23830
rect 23997 23810 24390 23824
rect 23997 23808 24003 23810
rect 23974 23805 24003 23808
rect 24387 23804 24390 23810
rect 24416 23804 24419 23830
rect 23652 23791 23681 23794
rect 23652 23774 23658 23791
rect 23675 23774 23681 23791
rect 23652 23771 23681 23774
rect 23744 23791 23773 23794
rect 23744 23774 23750 23791
rect 23767 23774 23773 23791
rect 23744 23771 23773 23774
rect 10955 23756 10958 23762
rect 9998 23742 10958 23756
rect 6916 23708 7850 23722
rect 9667 23702 9670 23728
rect 9696 23722 9699 23728
rect 9998 23722 10012 23742
rect 10955 23736 10958 23742
rect 10984 23756 10987 23762
rect 14635 23756 14638 23762
rect 10984 23742 14638 23756
rect 10984 23736 10987 23742
rect 14635 23736 14638 23742
rect 14664 23736 14667 23762
rect 9696 23708 10012 23722
rect 10059 23723 10088 23726
rect 9696 23702 9699 23708
rect 10059 23706 10065 23723
rect 10082 23722 10088 23723
rect 10219 23722 10222 23728
rect 10082 23708 10222 23722
rect 10082 23706 10088 23708
rect 10059 23703 10088 23706
rect 10219 23702 10222 23708
rect 10248 23702 10251 23728
rect 21306 23723 21335 23726
rect 21306 23706 21312 23723
rect 21329 23722 21335 23723
rect 21489 23722 21492 23728
rect 21329 23708 21492 23722
rect 21329 23706 21335 23708
rect 21306 23703 21335 23706
rect 21489 23702 21492 23708
rect 21518 23702 21521 23728
rect 23660 23722 23674 23771
rect 24525 23722 24528 23728
rect 23660 23708 24528 23722
rect 24525 23702 24528 23708
rect 24554 23722 24557 23728
rect 24664 23723 24693 23726
rect 24664 23722 24670 23723
rect 24554 23708 24670 23722
rect 24554 23702 24557 23708
rect 24664 23706 24670 23708
rect 24687 23706 24693 23723
rect 24664 23703 24693 23706
rect 3036 23640 29992 23688
rect 5067 23600 5070 23626
rect 5096 23620 5099 23626
rect 5251 23620 5254 23626
rect 5096 23606 5254 23620
rect 5096 23600 5099 23606
rect 5251 23600 5254 23606
rect 5280 23600 5283 23626
rect 5573 23600 5576 23626
rect 5602 23620 5605 23626
rect 6678 23621 6707 23624
rect 6678 23620 6684 23621
rect 5602 23606 6684 23620
rect 5602 23600 5605 23606
rect 6678 23604 6684 23606
rect 6701 23604 6707 23621
rect 12381 23620 12384 23626
rect 6678 23601 6707 23604
rect 8158 23606 12384 23620
rect 6401 23566 6404 23592
rect 6430 23566 6433 23592
rect 6033 23532 6036 23558
rect 6062 23552 6065 23558
rect 8158 23552 8172 23606
rect 6062 23538 8172 23552
rect 9484 23553 9513 23556
rect 6062 23532 6065 23538
rect 9484 23536 9490 23553
rect 9507 23552 9513 23553
rect 9507 23538 10196 23552
rect 9507 23536 9513 23538
rect 9484 23533 9513 23536
rect 3411 23498 3414 23524
rect 3440 23518 3443 23524
rect 5114 23519 5143 23522
rect 5114 23518 5120 23519
rect 3440 23504 5120 23518
rect 3440 23498 3443 23504
rect 5114 23502 5120 23504
rect 5137 23518 5143 23519
rect 5159 23518 5162 23524
rect 5137 23504 5162 23518
rect 5137 23502 5143 23504
rect 5114 23499 5143 23502
rect 5159 23498 5162 23504
rect 5188 23498 5191 23524
rect 5275 23519 5304 23522
rect 5275 23518 5281 23519
rect 5214 23504 5281 23518
rect 3457 23464 3460 23490
rect 3486 23484 3489 23490
rect 5214 23484 5228 23504
rect 5275 23502 5281 23504
rect 5298 23518 5304 23519
rect 5527 23518 5530 23524
rect 5298 23504 5530 23518
rect 5298 23502 5304 23504
rect 5275 23499 5304 23502
rect 5527 23498 5530 23504
rect 5556 23498 5559 23524
rect 6355 23498 6358 23524
rect 6384 23518 6387 23524
rect 6540 23519 6569 23522
rect 6540 23518 6546 23519
rect 6384 23504 6546 23518
rect 6384 23498 6387 23504
rect 6540 23502 6546 23504
rect 6563 23502 6569 23519
rect 6540 23499 6569 23502
rect 8149 23498 8152 23524
rect 8178 23498 8181 23524
rect 8287 23498 8290 23524
rect 8316 23522 8319 23524
rect 8316 23519 8334 23522
rect 8328 23502 8334 23519
rect 8885 23518 8888 23524
rect 8316 23499 8334 23502
rect 8388 23504 8888 23518
rect 8316 23498 8319 23499
rect 8388 23490 8402 23504
rect 8885 23498 8888 23504
rect 8914 23498 8917 23524
rect 9437 23498 9440 23524
rect 9466 23498 9469 23524
rect 9529 23498 9532 23524
rect 9558 23498 9561 23524
rect 10182 23522 10196 23538
rect 10174 23519 10203 23522
rect 10174 23502 10180 23519
rect 10197 23502 10203 23519
rect 10174 23499 10203 23502
rect 10219 23498 10222 23524
rect 10248 23498 10251 23524
rect 10274 23518 10288 23606
rect 12381 23600 12384 23606
rect 12410 23600 12413 23626
rect 18499 23600 18502 23626
rect 18528 23620 18531 23626
rect 20431 23624 20434 23626
rect 18546 23621 18575 23624
rect 18546 23620 18552 23621
rect 18528 23606 18552 23620
rect 18528 23600 18531 23606
rect 18546 23604 18552 23606
rect 18569 23604 18575 23621
rect 18546 23601 18575 23604
rect 20409 23621 20434 23624
rect 20409 23604 20415 23621
rect 20432 23604 20434 23621
rect 20409 23601 20434 23604
rect 20431 23600 20434 23601
rect 20460 23600 20463 23626
rect 17901 23566 17904 23592
rect 17930 23586 17933 23592
rect 17930 23572 18476 23586
rect 17930 23566 17933 23572
rect 10955 23532 10958 23558
rect 10984 23552 10987 23558
rect 10984 23538 11070 23552
rect 10984 23532 10987 23538
rect 10312 23519 10341 23522
rect 10312 23518 10318 23519
rect 10274 23504 10318 23518
rect 10312 23502 10318 23504
rect 10335 23502 10341 23519
rect 10312 23499 10341 23502
rect 10403 23498 10406 23524
rect 10432 23498 10435 23524
rect 11001 23498 11004 23524
rect 11030 23498 11033 23524
rect 11056 23518 11070 23538
rect 17073 23532 17076 23558
rect 17102 23552 17105 23558
rect 17856 23553 17885 23556
rect 17102 23538 17832 23552
rect 17102 23532 17105 23538
rect 11201 23519 11230 23522
rect 11201 23518 11207 23519
rect 11056 23504 11207 23518
rect 11201 23502 11207 23504
rect 11224 23502 11230 23519
rect 11415 23518 11418 23524
rect 11201 23499 11230 23502
rect 11332 23504 11418 23518
rect 5343 23488 5346 23490
rect 3486 23470 5228 23484
rect 5325 23485 5346 23488
rect 3486 23464 3489 23470
rect 5325 23468 5331 23485
rect 5325 23465 5346 23468
rect 5343 23464 5346 23465
rect 5372 23464 5375 23490
rect 8379 23488 8382 23490
rect 8361 23485 8382 23488
rect 8361 23468 8367 23485
rect 8361 23465 8382 23468
rect 8379 23464 8382 23465
rect 8408 23464 8411 23490
rect 10357 23464 10360 23490
rect 10386 23464 10389 23490
rect 11162 23485 11191 23488
rect 11162 23468 11168 23485
rect 11185 23484 11191 23485
rect 11332 23484 11346 23504
rect 11415 23498 11418 23504
rect 11444 23498 11447 23524
rect 12979 23498 12982 23524
rect 13008 23498 13011 23524
rect 13255 23498 13258 23524
rect 13284 23498 13287 23524
rect 16705 23498 16708 23524
rect 16734 23518 16737 23524
rect 17672 23519 17701 23522
rect 17672 23518 17678 23519
rect 16734 23504 17678 23518
rect 16734 23498 16737 23504
rect 17672 23502 17678 23504
rect 17695 23502 17701 23519
rect 17672 23499 17701 23502
rect 17764 23519 17793 23522
rect 17764 23502 17770 23519
rect 17787 23502 17793 23519
rect 17818 23518 17832 23538
rect 17856 23536 17862 23553
rect 17879 23552 17885 23553
rect 17947 23552 17950 23558
rect 17879 23538 17950 23552
rect 17879 23536 17885 23538
rect 17856 23533 17885 23536
rect 17947 23532 17950 23538
rect 17976 23552 17979 23558
rect 18131 23552 18134 23558
rect 17976 23538 18134 23552
rect 17976 23532 17979 23538
rect 18131 23532 18134 23538
rect 18160 23532 18163 23558
rect 18462 23556 18476 23572
rect 21213 23566 21216 23592
rect 21242 23566 21245 23592
rect 22685 23566 22688 23592
rect 22714 23586 22717 23592
rect 23605 23586 23608 23592
rect 22714 23572 23608 23586
rect 22714 23566 22717 23572
rect 23605 23566 23608 23572
rect 23634 23566 23637 23592
rect 18454 23553 18483 23556
rect 18454 23536 18460 23553
rect 18477 23536 18483 23553
rect 18454 23533 18483 23536
rect 18545 23532 18548 23558
rect 18574 23552 18577 23558
rect 18592 23553 18621 23556
rect 18592 23552 18598 23553
rect 18574 23538 18598 23552
rect 18574 23532 18577 23538
rect 18592 23536 18598 23538
rect 18615 23536 18621 23553
rect 18592 23533 18621 23536
rect 19373 23532 19376 23558
rect 19402 23532 19405 23558
rect 21397 23532 21400 23558
rect 21426 23552 21429 23558
rect 21719 23552 21722 23558
rect 21426 23538 21722 23552
rect 21426 23532 21429 23538
rect 21719 23532 21722 23538
rect 21748 23552 21751 23558
rect 21812 23553 21841 23556
rect 21812 23552 21818 23553
rect 21748 23538 21818 23552
rect 21748 23532 21751 23538
rect 21812 23536 21818 23538
rect 21835 23536 21841 23553
rect 21812 23533 21841 23536
rect 22847 23553 22876 23556
rect 22847 23536 22853 23553
rect 22870 23552 22876 23553
rect 23146 23553 23175 23556
rect 23146 23552 23152 23553
rect 22870 23538 23152 23552
rect 22870 23536 22876 23538
rect 22847 23533 22876 23536
rect 23146 23536 23152 23538
rect 23169 23536 23175 23553
rect 23146 23533 23175 23536
rect 17902 23519 17931 23522
rect 17902 23518 17908 23519
rect 17818 23504 17908 23518
rect 17764 23499 17793 23502
rect 17902 23502 17908 23504
rect 17925 23502 17931 23519
rect 17902 23499 17931 23502
rect 18500 23519 18529 23522
rect 18500 23502 18506 23519
rect 18523 23502 18529 23519
rect 18500 23499 18529 23502
rect 19535 23519 19564 23522
rect 19535 23502 19541 23519
rect 19558 23518 19564 23519
rect 20017 23518 20020 23524
rect 19558 23504 20020 23518
rect 19558 23502 19564 23504
rect 19535 23499 19564 23502
rect 11185 23470 11346 23484
rect 11185 23468 11191 23470
rect 11162 23465 11191 23468
rect 17257 23464 17260 23490
rect 17286 23484 17289 23490
rect 17772 23484 17786 23499
rect 17809 23484 17812 23490
rect 17286 23470 17812 23484
rect 17286 23464 17289 23470
rect 17809 23464 17812 23470
rect 17838 23464 17841 23490
rect 18508 23484 18522 23499
rect 20017 23498 20020 23504
rect 20046 23498 20049 23524
rect 21351 23498 21354 23524
rect 21380 23498 21383 23524
rect 21949 23498 21952 23524
rect 21978 23522 21981 23524
rect 21978 23519 22002 23522
rect 21978 23502 21979 23519
rect 21996 23518 22002 23519
rect 23192 23519 23221 23522
rect 23192 23518 23198 23519
rect 21996 23504 23198 23518
rect 21996 23502 22002 23504
rect 21978 23499 22002 23502
rect 23192 23502 23198 23504
rect 23215 23518 23221 23519
rect 23421 23518 23424 23524
rect 23215 23504 23424 23518
rect 23215 23502 23221 23504
rect 23192 23499 23221 23502
rect 21978 23498 21981 23499
rect 23421 23498 23424 23504
rect 23450 23498 23453 23524
rect 24433 23522 24436 23524
rect 24296 23519 24325 23522
rect 24296 23502 24302 23519
rect 24319 23502 24325 23519
rect 24430 23518 24436 23522
rect 24413 23504 24436 23518
rect 24296 23499 24325 23502
rect 24430 23499 24436 23504
rect 18591 23484 18594 23490
rect 18508 23470 18594 23484
rect 18591 23464 18594 23470
rect 18620 23464 18623 23490
rect 19419 23464 19422 23490
rect 19448 23484 19451 23490
rect 19581 23485 19610 23488
rect 19581 23484 19587 23485
rect 19448 23470 19587 23484
rect 19448 23464 19451 23470
rect 19581 23468 19587 23470
rect 19604 23468 19610 23485
rect 19581 23465 19610 23468
rect 21214 23485 21243 23488
rect 21214 23468 21220 23485
rect 21237 23484 21243 23485
rect 21259 23484 21262 23490
rect 21237 23470 21262 23484
rect 21237 23468 21243 23470
rect 21214 23465 21243 23468
rect 21259 23464 21262 23470
rect 21288 23464 21291 23490
rect 22041 23488 22044 23490
rect 22023 23485 22044 23488
rect 22023 23468 22029 23485
rect 22023 23465 22044 23468
rect 22041 23464 22044 23465
rect 22070 23464 22073 23490
rect 24304 23484 24318 23499
rect 24433 23498 24436 23499
rect 24462 23498 24465 23524
rect 24387 23484 24390 23490
rect 24304 23470 24390 23484
rect 24387 23464 24390 23470
rect 24416 23464 24419 23490
rect 6149 23451 6178 23454
rect 6149 23434 6155 23451
rect 6172 23450 6178 23451
rect 6263 23450 6266 23456
rect 6172 23436 6266 23450
rect 6172 23434 6178 23436
rect 6149 23431 6178 23434
rect 6263 23430 6266 23436
rect 6292 23430 6295 23456
rect 6309 23430 6312 23456
rect 6338 23450 6341 23456
rect 6494 23451 6523 23454
rect 6494 23450 6500 23451
rect 6338 23436 6500 23450
rect 6338 23430 6341 23436
rect 6494 23434 6500 23436
rect 6517 23434 6523 23451
rect 6494 23431 6523 23434
rect 6586 23451 6615 23454
rect 6586 23434 6592 23451
rect 6609 23450 6615 23451
rect 8195 23450 8198 23456
rect 6609 23436 8198 23450
rect 6609 23434 6615 23436
rect 6586 23431 6615 23434
rect 8195 23430 8198 23436
rect 8224 23430 8227 23456
rect 9185 23451 9214 23454
rect 9185 23434 9191 23451
rect 9208 23450 9214 23451
rect 9391 23450 9394 23456
rect 9208 23436 9394 23450
rect 9208 23434 9214 23436
rect 9185 23431 9214 23434
rect 9391 23430 9394 23436
rect 9420 23430 9423 23456
rect 10266 23451 10295 23454
rect 10266 23434 10272 23451
rect 10289 23450 10295 23451
rect 10633 23450 10636 23456
rect 10289 23436 10636 23450
rect 10289 23434 10295 23436
rect 10266 23431 10295 23434
rect 10633 23430 10636 23436
rect 10662 23430 10665 23456
rect 12013 23430 12016 23456
rect 12042 23454 12045 23456
rect 12042 23451 12066 23454
rect 12042 23434 12043 23451
rect 12060 23434 12066 23451
rect 12042 23431 12066 23434
rect 12042 23430 12045 23431
rect 12887 23430 12890 23456
rect 12916 23450 12919 23456
rect 13026 23451 13055 23454
rect 13026 23450 13032 23451
rect 12916 23436 13032 23450
rect 12916 23430 12919 23436
rect 13026 23434 13032 23436
rect 13049 23434 13055 23451
rect 13026 23431 13055 23434
rect 15233 23430 15236 23456
rect 15262 23450 15265 23456
rect 15831 23450 15834 23456
rect 15262 23436 15834 23450
rect 15262 23430 15265 23436
rect 15831 23430 15834 23436
rect 15860 23450 15863 23456
rect 17947 23450 17950 23456
rect 15860 23436 17950 23450
rect 15860 23430 15863 23436
rect 17947 23430 17950 23436
rect 17976 23430 17979 23456
rect 21306 23451 21335 23454
rect 21306 23434 21312 23451
rect 21329 23450 21335 23451
rect 21581 23450 21584 23456
rect 21329 23436 21584 23450
rect 21329 23434 21335 23436
rect 21306 23431 21335 23434
rect 21581 23430 21584 23436
rect 21610 23430 21613 23456
rect 23375 23430 23378 23456
rect 23404 23430 23407 23456
rect 24801 23430 24804 23456
rect 24830 23450 24833 23456
rect 24986 23451 25015 23454
rect 24986 23450 24992 23451
rect 24830 23436 24992 23450
rect 24830 23430 24833 23436
rect 24986 23434 24992 23436
rect 25009 23434 25015 23451
rect 24986 23431 25015 23434
rect 3036 23368 29992 23416
rect 10243 23349 10272 23352
rect 10243 23332 10249 23349
rect 10266 23348 10272 23349
rect 10357 23348 10360 23354
rect 10266 23334 10360 23348
rect 10266 23332 10272 23334
rect 10243 23329 10272 23332
rect 10357 23328 10360 23334
rect 10386 23328 10389 23354
rect 10679 23328 10682 23354
rect 10708 23328 10711 23354
rect 10725 23328 10728 23354
rect 10754 23328 10757 23354
rect 10817 23328 10820 23354
rect 10846 23328 10849 23354
rect 11033 23334 12266 23348
rect 6263 23294 6266 23320
rect 6292 23294 6295 23320
rect 6356 23315 6385 23318
rect 6356 23298 6362 23315
rect 6379 23314 6385 23315
rect 6631 23314 6634 23320
rect 6379 23300 6634 23314
rect 6379 23298 6385 23300
rect 6356 23295 6385 23298
rect 6631 23294 6634 23300
rect 6660 23294 6663 23320
rect 9253 23294 9256 23320
rect 9282 23314 9285 23320
rect 9415 23315 9444 23318
rect 9415 23314 9421 23315
rect 9282 23300 9421 23314
rect 9282 23294 9285 23300
rect 9415 23298 9421 23300
rect 9438 23298 9444 23315
rect 9415 23295 9444 23298
rect 10403 23294 10406 23320
rect 10432 23314 10435 23320
rect 11033 23314 11047 23334
rect 10432 23300 11047 23314
rect 11562 23300 11714 23314
rect 10432 23294 10435 23300
rect 6401 23260 6404 23286
rect 6430 23260 6433 23286
rect 6466 23281 6495 23284
rect 6466 23264 6472 23281
rect 6489 23280 6495 23281
rect 6723 23280 6726 23286
rect 6489 23266 6726 23280
rect 6489 23264 6495 23266
rect 6466 23261 6495 23264
rect 6723 23260 6726 23266
rect 6752 23260 6755 23286
rect 9161 23260 9164 23286
rect 9190 23280 9193 23286
rect 9345 23280 9348 23286
rect 9374 23284 9377 23286
rect 9374 23281 9392 23284
rect 9190 23266 9348 23280
rect 9190 23260 9193 23266
rect 9345 23260 9348 23266
rect 9386 23264 9392 23281
rect 9374 23261 9392 23264
rect 9374 23260 9377 23261
rect 10633 23260 10636 23286
rect 10662 23260 10665 23286
rect 10863 23260 10866 23286
rect 10892 23280 10895 23286
rect 11562 23284 11576 23300
rect 11554 23281 11583 23284
rect 11554 23280 11560 23281
rect 10892 23266 11560 23280
rect 10892 23260 10895 23266
rect 11554 23264 11560 23266
rect 11577 23264 11583 23281
rect 11554 23261 11583 23264
rect 11645 23260 11648 23286
rect 11674 23260 11677 23286
rect 6309 23226 6312 23252
rect 6338 23226 6341 23252
rect 9023 23226 9026 23252
rect 9052 23246 9055 23252
rect 9208 23247 9237 23250
rect 9208 23246 9214 23247
rect 9052 23232 9214 23246
rect 9052 23226 9055 23232
rect 9208 23230 9214 23232
rect 9231 23230 9237 23247
rect 9208 23227 9237 23230
rect 10818 23247 10847 23250
rect 10818 23230 10824 23247
rect 10841 23246 10847 23247
rect 11600 23247 11629 23250
rect 11600 23246 11606 23247
rect 10841 23232 11606 23246
rect 10841 23230 10847 23232
rect 10818 23227 10847 23230
rect 11600 23230 11606 23232
rect 11623 23230 11629 23247
rect 11600 23227 11629 23230
rect 11700 23212 11714 23300
rect 12013 23294 12016 23320
rect 12042 23294 12045 23320
rect 12105 23294 12108 23320
rect 12134 23294 12137 23320
rect 12252 23314 12266 23334
rect 14635 23328 14638 23354
rect 14664 23328 14667 23354
rect 15233 23348 15236 23354
rect 14690 23334 15236 23348
rect 14690 23314 14704 23334
rect 15233 23328 15236 23334
rect 15262 23328 15265 23354
rect 17119 23328 17122 23354
rect 17148 23328 17151 23354
rect 17947 23328 17950 23354
rect 17976 23328 17979 23354
rect 14957 23314 14960 23320
rect 12252 23300 14704 23314
rect 14736 23300 14960 23314
rect 12151 23260 12154 23286
rect 12180 23260 12183 23286
rect 12208 23281 12237 23284
rect 12208 23264 12214 23281
rect 12231 23280 12237 23281
rect 12252 23280 12266 23300
rect 12231 23266 12266 23280
rect 12231 23264 12237 23266
rect 12208 23261 12237 23264
rect 13117 23260 13120 23286
rect 13146 23260 13149 23286
rect 13255 23260 13258 23286
rect 13284 23280 13287 23286
rect 14736 23284 14750 23300
rect 14957 23294 14960 23300
rect 14986 23294 14989 23320
rect 17257 23314 17260 23320
rect 17128 23300 17260 23314
rect 14728 23281 14757 23284
rect 13284 23266 14244 23280
rect 13284 23260 13287 23266
rect 12060 23247 12089 23250
rect 12060 23230 12066 23247
rect 12083 23246 12089 23247
rect 12289 23246 12292 23252
rect 12083 23232 12292 23246
rect 12083 23230 12089 23232
rect 12060 23227 12089 23230
rect 12289 23226 12292 23232
rect 12318 23226 12321 23252
rect 12841 23226 12844 23252
rect 12870 23246 12873 23252
rect 13210 23247 13239 23250
rect 13210 23246 13216 23247
rect 12870 23232 13216 23246
rect 12870 23226 12873 23232
rect 13210 23230 13216 23232
rect 13233 23230 13239 23247
rect 14230 23246 14244 23266
rect 14728 23264 14734 23281
rect 14751 23264 14757 23281
rect 14728 23261 14757 23264
rect 14866 23281 14895 23284
rect 14866 23264 14872 23281
rect 14889 23280 14895 23281
rect 14911 23280 14914 23286
rect 14889 23266 14914 23280
rect 14889 23264 14895 23266
rect 14866 23261 14895 23264
rect 14874 23246 14888 23261
rect 14911 23260 14914 23266
rect 14940 23260 14943 23286
rect 16291 23260 16294 23286
rect 16320 23260 16323 23286
rect 16521 23260 16524 23286
rect 16550 23280 16553 23286
rect 17128 23284 17142 23300
rect 17257 23294 17260 23300
rect 17286 23294 17289 23320
rect 20566 23315 20595 23318
rect 19290 23300 20546 23314
rect 17120 23281 17149 23284
rect 16550 23266 16682 23280
rect 16550 23260 16553 23266
rect 14230 23232 14888 23246
rect 14958 23247 14987 23250
rect 13210 23227 13239 23230
rect 14958 23230 14964 23247
rect 14981 23246 14987 23247
rect 15003 23246 15006 23252
rect 14981 23232 15006 23246
rect 14981 23230 14987 23232
rect 14958 23227 14987 23230
rect 15003 23226 15006 23232
rect 15032 23226 15035 23252
rect 16567 23226 16570 23252
rect 16596 23226 16599 23252
rect 16668 23246 16682 23266
rect 17120 23264 17126 23281
rect 17143 23264 17149 23281
rect 17120 23261 17149 23264
rect 17165 23260 17168 23286
rect 17194 23280 17197 23286
rect 17212 23281 17241 23284
rect 17212 23280 17218 23281
rect 17194 23266 17218 23280
rect 17194 23260 17197 23266
rect 17212 23264 17218 23266
rect 17235 23264 17241 23281
rect 17212 23261 17241 23264
rect 17901 23260 17904 23286
rect 17930 23260 17933 23286
rect 18131 23260 18134 23286
rect 18160 23260 18163 23286
rect 18499 23260 18502 23286
rect 18528 23280 18531 23286
rect 19290 23284 19304 23300
rect 19006 23281 19035 23284
rect 19006 23280 19012 23281
rect 18528 23266 19012 23280
rect 18528 23260 18531 23266
rect 19006 23264 19012 23266
rect 19029 23264 19035 23281
rect 19006 23261 19035 23264
rect 19282 23281 19311 23284
rect 19282 23264 19288 23281
rect 19305 23264 19311 23281
rect 19282 23261 19311 23264
rect 19374 23281 19403 23284
rect 19374 23264 19380 23281
rect 19397 23280 19403 23281
rect 19419 23280 19422 23286
rect 19397 23266 19422 23280
rect 19397 23264 19403 23266
rect 19374 23261 19403 23264
rect 19419 23260 19422 23266
rect 19448 23260 19451 23286
rect 20532 23280 20546 23300
rect 20566 23298 20572 23315
rect 20589 23314 20595 23315
rect 21213 23314 21216 23320
rect 20589 23300 21216 23314
rect 20589 23298 20595 23300
rect 20566 23295 20595 23298
rect 21213 23294 21216 23300
rect 21242 23294 21245 23320
rect 21489 23318 21492 23320
rect 21486 23314 21492 23318
rect 21469 23300 21492 23314
rect 21486 23295 21492 23300
rect 21489 23294 21492 23295
rect 21518 23294 21521 23320
rect 21075 23280 21078 23286
rect 20532 23266 21078 23280
rect 21075 23260 21078 23266
rect 21104 23260 21107 23286
rect 21351 23260 21354 23286
rect 21380 23260 21383 23286
rect 17304 23247 17333 23250
rect 17304 23246 17310 23247
rect 16668 23232 17310 23246
rect 17304 23230 17310 23232
rect 17327 23230 17333 23247
rect 20432 23247 20461 23250
rect 20432 23246 20438 23247
rect 17304 23227 17333 23230
rect 19382 23232 20438 23246
rect 19382 23218 19396 23232
rect 20432 23230 20438 23232
rect 20455 23230 20461 23247
rect 20432 23227 20461 23230
rect 16153 23212 16156 23218
rect 11700 23198 16156 23212
rect 16153 23192 16156 23198
rect 16182 23192 16185 23218
rect 19373 23192 19376 23218
rect 19402 23192 19405 23218
rect 6723 23158 6726 23184
rect 6752 23178 6755 23184
rect 10403 23178 10406 23184
rect 6752 23164 10406 23178
rect 6752 23158 6755 23164
rect 10403 23158 10406 23164
rect 10432 23158 10435 23184
rect 12105 23158 12108 23184
rect 12134 23178 12137 23184
rect 15233 23178 15236 23184
rect 12134 23164 15236 23178
rect 12134 23158 12137 23164
rect 15233 23158 15236 23164
rect 15262 23158 15265 23184
rect 20440 23178 20454 23227
rect 21360 23212 21374 23260
rect 21084 23198 21374 23212
rect 21084 23178 21098 23198
rect 20440 23164 21098 23178
rect 21121 23158 21124 23184
rect 21150 23158 21153 23184
rect 22041 23158 22044 23184
rect 22070 23158 22073 23184
rect 3036 23096 29992 23144
rect 6447 23056 6450 23082
rect 6476 23076 6479 23082
rect 6517 23077 6546 23080
rect 6517 23076 6523 23077
rect 6476 23062 6523 23076
rect 6476 23056 6479 23062
rect 6517 23060 6523 23062
rect 6540 23060 6546 23077
rect 6517 23057 6546 23060
rect 9346 23077 9375 23080
rect 9346 23060 9352 23077
rect 9369 23076 9375 23077
rect 9529 23076 9532 23082
rect 9369 23062 9532 23076
rect 9369 23060 9375 23062
rect 9346 23057 9375 23060
rect 9529 23056 9532 23062
rect 9558 23056 9561 23082
rect 12151 23080 12154 23082
rect 12129 23077 12154 23080
rect 11102 23062 12082 23076
rect 6631 23022 6634 23048
rect 6660 23042 6663 23048
rect 10863 23042 10866 23048
rect 6660 23028 10866 23042
rect 6660 23022 6663 23028
rect 10863 23022 10866 23028
rect 10892 23022 10895 23048
rect 4837 22988 4840 23014
rect 4866 23008 4869 23014
rect 4866 22994 5550 23008
rect 4866 22988 4869 22994
rect 5159 22954 5162 22980
rect 5188 22974 5191 22980
rect 5297 22974 5300 22980
rect 5188 22960 5300 22974
rect 5188 22954 5191 22960
rect 5297 22954 5300 22960
rect 5326 22974 5329 22980
rect 5482 22975 5511 22978
rect 5482 22974 5488 22975
rect 5326 22960 5488 22974
rect 5326 22954 5329 22960
rect 5482 22958 5488 22960
rect 5505 22958 5511 22975
rect 5536 22974 5550 22994
rect 9253 22988 9256 23014
rect 9282 23008 9285 23014
rect 11102 23008 11116 23062
rect 12068 23008 12082 23062
rect 12129 23060 12135 23077
rect 12152 23060 12154 23077
rect 12129 23057 12154 23060
rect 12151 23056 12154 23057
rect 12180 23056 12183 23082
rect 16521 23056 16524 23082
rect 16550 23076 16553 23082
rect 16660 23077 16689 23080
rect 16660 23076 16666 23077
rect 16550 23062 16666 23076
rect 16550 23056 16553 23062
rect 16660 23060 16666 23062
rect 16683 23060 16689 23077
rect 16660 23057 16689 23060
rect 17533 23056 17536 23082
rect 17562 23056 17565 23082
rect 21259 23056 21262 23082
rect 21288 23076 21291 23082
rect 21306 23077 21335 23080
rect 21306 23076 21312 23077
rect 21288 23062 21312 23076
rect 21288 23056 21291 23062
rect 21306 23060 21312 23062
rect 21329 23060 21335 23077
rect 21306 23057 21335 23060
rect 21673 23056 21676 23082
rect 21702 23056 21705 23082
rect 22685 23056 22688 23082
rect 22714 23056 22717 23082
rect 14221 23022 14224 23048
rect 14250 23042 14253 23048
rect 18407 23042 18410 23048
rect 14250 23028 18410 23042
rect 14250 23022 14253 23028
rect 18407 23022 18410 23028
rect 18436 23042 18439 23048
rect 18499 23042 18502 23048
rect 18436 23028 18502 23042
rect 18436 23022 18439 23028
rect 18499 23022 18502 23028
rect 18528 23022 18531 23048
rect 19880 23043 19909 23046
rect 19880 23026 19886 23043
rect 19903 23026 19909 23043
rect 19880 23023 19909 23026
rect 14681 23008 14684 23014
rect 9282 22994 11162 23008
rect 12068 22994 14684 23008
rect 9282 22988 9285 22994
rect 9300 22975 9329 22978
rect 9300 22974 9306 22975
rect 5536 22960 9306 22974
rect 5482 22955 5511 22958
rect 9300 22958 9306 22960
rect 9323 22958 9329 22975
rect 9300 22955 9329 22958
rect 5251 22920 5254 22946
rect 5280 22940 5283 22946
rect 5435 22940 5438 22946
rect 5280 22926 5438 22940
rect 5280 22920 5283 22926
rect 5435 22920 5438 22926
rect 5464 22920 5467 22946
rect 5527 22920 5530 22946
rect 5556 22940 5559 22946
rect 5642 22941 5671 22944
rect 5642 22940 5648 22941
rect 5556 22926 5648 22940
rect 5556 22920 5559 22926
rect 5642 22924 5648 22926
rect 5665 22924 5671 22941
rect 5642 22921 5671 22924
rect 5693 22941 5722 22944
rect 5693 22924 5699 22941
rect 5716 22940 5722 22941
rect 5757 22940 5760 22946
rect 5716 22926 5760 22940
rect 5716 22924 5722 22926
rect 5693 22921 5722 22924
rect 5757 22920 5760 22926
rect 5786 22920 5789 22946
rect 9308 22940 9322 22955
rect 9391 22954 9394 22980
rect 9420 22954 9423 22980
rect 11047 22954 11050 22980
rect 11076 22974 11079 22980
rect 11094 22975 11123 22978
rect 11094 22974 11100 22975
rect 11076 22960 11100 22974
rect 11076 22954 11079 22960
rect 11094 22958 11100 22960
rect 11117 22958 11123 22975
rect 11094 22955 11123 22958
rect 10265 22940 10268 22946
rect 9308 22926 10268 22940
rect 10265 22920 10268 22926
rect 10294 22920 10297 22946
rect 11148 22940 11162 22994
rect 14681 22988 14684 22994
rect 14710 22988 14713 23014
rect 15095 22988 15098 23014
rect 15124 22988 15127 23014
rect 17671 22988 17674 23014
rect 17700 23008 17703 23014
rect 17856 23009 17885 23012
rect 17856 23008 17862 23009
rect 17700 22994 17862 23008
rect 17700 22988 17703 22994
rect 17856 22992 17862 22994
rect 17879 22992 17885 23009
rect 17856 22989 17885 22992
rect 17948 23009 17977 23012
rect 17948 22992 17954 23009
rect 17971 23008 17977 23009
rect 18545 23008 18548 23014
rect 17971 22994 18548 23008
rect 17971 22992 17977 22994
rect 17948 22989 17977 22992
rect 18545 22988 18548 22994
rect 18574 22988 18577 23014
rect 19649 22988 19652 23014
rect 19678 22988 19681 23014
rect 19888 23008 19902 23023
rect 21075 23022 21078 23048
rect 21104 23042 21107 23048
rect 21104 23028 22478 23042
rect 21104 23022 21107 23028
rect 20202 23009 20231 23012
rect 20202 23008 20208 23009
rect 19888 22994 20208 23008
rect 20202 22992 20208 22994
rect 20225 22992 20231 23009
rect 20202 22989 20231 22992
rect 21213 22988 21216 23014
rect 21242 22988 21245 23014
rect 21305 22988 21308 23014
rect 21334 23008 21337 23014
rect 21352 23009 21381 23012
rect 21352 23008 21358 23009
rect 21334 22994 21358 23008
rect 21334 22988 21337 22994
rect 21352 22992 21358 22994
rect 21375 23008 21381 23009
rect 21720 23009 21749 23012
rect 21720 23008 21726 23009
rect 21375 22994 21726 23008
rect 21375 22992 21381 22994
rect 21352 22989 21381 22992
rect 21720 22992 21726 22994
rect 21743 22992 21749 23009
rect 21720 22989 21749 22992
rect 22464 23008 22478 23028
rect 22464 22994 23076 23008
rect 11255 22975 11284 22978
rect 11255 22958 11261 22975
rect 11278 22974 11284 22975
rect 11415 22974 11418 22980
rect 11278 22960 11418 22974
rect 11278 22958 11284 22960
rect 11255 22955 11284 22958
rect 11415 22954 11418 22960
rect 11444 22954 11447 22980
rect 13117 22954 13120 22980
rect 13146 22974 13149 22980
rect 13348 22975 13377 22978
rect 13348 22974 13354 22975
rect 13146 22960 13354 22974
rect 13146 22954 13149 22960
rect 13348 22958 13354 22960
rect 13371 22974 13377 22975
rect 13393 22974 13396 22980
rect 13371 22960 13396 22974
rect 13371 22958 13377 22960
rect 13348 22955 13377 22958
rect 13393 22954 13396 22960
rect 13422 22954 13425 22980
rect 13624 22975 13653 22978
rect 13624 22958 13630 22975
rect 13647 22974 13653 22975
rect 14497 22974 14500 22980
rect 13647 22960 14500 22974
rect 13647 22958 13653 22960
rect 13624 22955 13653 22958
rect 14497 22954 14500 22960
rect 14526 22954 14529 22980
rect 14957 22954 14960 22980
rect 14986 22954 14989 22980
rect 15050 22975 15079 22978
rect 15050 22958 15056 22975
rect 15073 22958 15079 22975
rect 15050 22955 15079 22958
rect 16108 22975 16137 22978
rect 16108 22958 16114 22975
rect 16131 22958 16137 22975
rect 16108 22955 16137 22958
rect 11301 22941 11330 22944
rect 11301 22940 11307 22941
rect 11148 22926 11307 22940
rect 11301 22924 11307 22926
rect 11324 22924 11330 22941
rect 11301 22921 11330 22924
rect 13716 22941 13745 22944
rect 13716 22924 13722 22941
rect 13739 22940 13745 22941
rect 14405 22940 14408 22946
rect 13739 22926 14408 22940
rect 13739 22924 13745 22926
rect 13716 22921 13745 22924
rect 14405 22920 14408 22926
rect 14434 22920 14437 22946
rect 14506 22940 14520 22954
rect 15058 22940 15072 22955
rect 14506 22926 15072 22940
rect 16116 22940 16130 22955
rect 16245 22954 16248 22980
rect 16274 22974 16277 22980
rect 16521 22974 16524 22980
rect 16274 22960 16524 22974
rect 16274 22954 16277 22960
rect 16521 22954 16524 22960
rect 16550 22954 16553 22980
rect 16660 22975 16689 22978
rect 16660 22958 16666 22975
rect 16683 22958 16689 22975
rect 16660 22955 16689 22958
rect 16429 22940 16432 22946
rect 16116 22926 16432 22940
rect 16429 22920 16432 22926
rect 16458 22920 16461 22946
rect 16668 22940 16682 22955
rect 16705 22954 16708 22980
rect 16734 22974 16737 22980
rect 16890 22975 16919 22978
rect 16890 22974 16896 22975
rect 16734 22960 16896 22974
rect 16734 22954 16737 22960
rect 16890 22958 16896 22960
rect 16913 22958 16919 22975
rect 16890 22955 16919 22958
rect 17487 22954 17490 22980
rect 17516 22954 17519 22980
rect 17579 22954 17582 22980
rect 17608 22954 17611 22980
rect 17809 22954 17812 22980
rect 17838 22954 17841 22980
rect 19696 22975 19725 22978
rect 19696 22958 19702 22975
rect 19719 22974 19725 22975
rect 20155 22974 20158 22980
rect 19719 22960 20158 22974
rect 19719 22958 19725 22960
rect 19696 22955 19725 22958
rect 20155 22954 20158 22960
rect 20184 22954 20187 22980
rect 20339 22954 20342 22980
rect 20368 22954 20371 22980
rect 21121 22974 21124 22980
rect 20693 22960 21124 22974
rect 17395 22940 17398 22946
rect 16668 22926 17398 22940
rect 17395 22920 17398 22926
rect 17424 22940 17427 22946
rect 17901 22940 17904 22946
rect 17424 22926 17904 22940
rect 17424 22920 17427 22926
rect 17901 22920 17904 22926
rect 17930 22920 17933 22946
rect 19787 22920 19790 22946
rect 19816 22940 19819 22946
rect 20693 22940 20707 22960
rect 21121 22954 21124 22960
rect 21150 22974 21153 22980
rect 21260 22975 21289 22978
rect 21260 22974 21266 22975
rect 21150 22960 21266 22974
rect 21150 22954 21153 22960
rect 21260 22958 21266 22960
rect 21283 22958 21289 22975
rect 21260 22955 21289 22958
rect 21581 22954 21584 22980
rect 21610 22954 21613 22980
rect 21627 22954 21630 22980
rect 21656 22974 21659 22980
rect 22041 22974 22044 22980
rect 21656 22960 22044 22974
rect 21656 22954 21659 22960
rect 22041 22954 22044 22960
rect 22070 22954 22073 22980
rect 22464 22978 22478 22994
rect 22456 22975 22485 22978
rect 22456 22958 22462 22975
rect 22479 22958 22485 22975
rect 22456 22955 22485 22958
rect 22823 22954 22826 22980
rect 22852 22974 22855 22980
rect 23062 22978 23076 22994
rect 22962 22975 22991 22978
rect 22962 22974 22968 22975
rect 22852 22960 22968 22974
rect 22852 22954 22855 22960
rect 22962 22958 22968 22960
rect 22985 22958 22991 22975
rect 22962 22955 22991 22958
rect 23054 22975 23083 22978
rect 23054 22958 23060 22975
rect 23077 22974 23083 22975
rect 23191 22974 23194 22980
rect 23077 22960 23194 22974
rect 23077 22958 23083 22960
rect 23054 22955 23083 22958
rect 23191 22954 23194 22960
rect 23220 22954 23223 22980
rect 24387 22954 24390 22980
rect 24416 22974 24419 22980
rect 24618 22975 24647 22978
rect 24618 22974 24624 22975
rect 24416 22960 24624 22974
rect 24416 22954 24419 22960
rect 24618 22958 24624 22960
rect 24641 22958 24647 22975
rect 24618 22955 24647 22958
rect 19816 22926 20707 22940
rect 21590 22940 21604 22954
rect 22732 22941 22761 22944
rect 22732 22940 22738 22941
rect 21590 22926 22738 22940
rect 19816 22920 19819 22926
rect 5941 22886 5944 22912
rect 5970 22906 5973 22912
rect 9253 22906 9256 22912
rect 5970 22892 9256 22906
rect 5970 22886 5973 22892
rect 9253 22886 9256 22892
rect 9282 22886 9285 22912
rect 11553 22886 11556 22912
rect 11582 22906 11585 22912
rect 13394 22907 13423 22910
rect 13394 22906 13400 22907
rect 11582 22892 13400 22906
rect 11582 22886 11585 22892
rect 13394 22890 13400 22892
rect 13417 22890 13423 22907
rect 13394 22887 13423 22890
rect 16108 22907 16137 22910
rect 16108 22890 16114 22907
rect 16131 22906 16137 22907
rect 16153 22906 16156 22912
rect 16131 22892 16156 22906
rect 16131 22890 16137 22892
rect 16108 22887 16137 22890
rect 16153 22886 16156 22892
rect 16182 22886 16185 22912
rect 17947 22886 17950 22912
rect 17976 22886 17979 22912
rect 20662 22907 20691 22910
rect 20662 22890 20668 22907
rect 20685 22906 20691 22907
rect 20845 22906 20848 22912
rect 20685 22892 20848 22906
rect 20685 22890 20691 22892
rect 20662 22887 20691 22890
rect 20845 22886 20848 22892
rect 20874 22886 20877 22912
rect 21213 22886 21216 22912
rect 21242 22906 21245 22912
rect 21590 22906 21604 22926
rect 22732 22924 22738 22926
rect 22755 22924 22761 22941
rect 22732 22921 22761 22924
rect 24525 22920 24528 22946
rect 24554 22940 24557 22946
rect 24847 22944 24850 22946
rect 24778 22941 24807 22944
rect 24778 22940 24784 22941
rect 24554 22926 24784 22940
rect 24554 22920 24557 22926
rect 24778 22924 24784 22926
rect 24801 22924 24807 22941
rect 24778 22921 24807 22924
rect 24829 22941 24850 22944
rect 24829 22924 24835 22941
rect 24829 22921 24850 22924
rect 24847 22920 24850 22921
rect 24876 22920 24879 22946
rect 21242 22892 21604 22906
rect 23008 22907 23037 22910
rect 21242 22886 21245 22892
rect 23008 22890 23014 22907
rect 23031 22906 23037 22907
rect 23375 22906 23378 22912
rect 23031 22892 23378 22906
rect 23031 22890 23037 22892
rect 23008 22887 23037 22890
rect 23375 22886 23378 22892
rect 23404 22886 23407 22912
rect 25629 22886 25632 22912
rect 25658 22910 25661 22912
rect 25658 22907 25682 22910
rect 25658 22890 25659 22907
rect 25676 22890 25682 22907
rect 25658 22887 25682 22890
rect 25658 22886 25661 22887
rect 3036 22824 29992 22872
rect 11071 22805 11100 22808
rect 11071 22788 11077 22805
rect 11094 22804 11100 22805
rect 11645 22804 11648 22810
rect 11094 22790 11648 22804
rect 11094 22788 11100 22790
rect 11071 22785 11100 22788
rect 11645 22784 11648 22790
rect 11674 22784 11677 22810
rect 14543 22784 14546 22810
rect 14572 22804 14575 22810
rect 14681 22804 14684 22810
rect 14572 22790 14684 22804
rect 14572 22784 14575 22790
rect 14681 22784 14684 22790
rect 14710 22784 14713 22810
rect 14957 22784 14960 22810
rect 14986 22784 14989 22810
rect 18316 22805 18345 22808
rect 18316 22788 18322 22805
rect 18339 22788 18345 22805
rect 18316 22785 18345 22788
rect 19374 22805 19403 22808
rect 19374 22788 19380 22805
rect 19397 22804 19403 22805
rect 19649 22804 19652 22810
rect 19397 22790 19652 22804
rect 19397 22788 19403 22790
rect 19374 22785 19403 22788
rect 9713 22750 9716 22776
rect 9742 22770 9745 22776
rect 14966 22770 14980 22784
rect 17487 22770 17490 22776
rect 9742 22756 10265 22770
rect 9742 22750 9745 22756
rect 3549 22716 3552 22742
rect 3578 22740 3581 22742
rect 3578 22737 3596 22740
rect 3590 22720 3596 22737
rect 3578 22717 3596 22720
rect 3611 22737 3640 22740
rect 3611 22720 3617 22737
rect 3634 22736 3640 22737
rect 3687 22736 3690 22742
rect 3634 22722 3690 22736
rect 3634 22720 3640 22722
rect 3611 22717 3640 22720
rect 3578 22716 3581 22717
rect 3687 22716 3690 22722
rect 3716 22716 3719 22742
rect 7321 22716 7324 22742
rect 7350 22736 7353 22742
rect 7431 22737 7460 22740
rect 7431 22736 7437 22737
rect 7350 22722 7437 22736
rect 7350 22716 7353 22722
rect 7431 22720 7437 22722
rect 7454 22720 7460 22737
rect 7431 22717 7460 22720
rect 7475 22737 7504 22740
rect 7475 22720 7481 22737
rect 7498 22736 7504 22737
rect 7551 22736 7554 22742
rect 7498 22722 7554 22736
rect 7498 22720 7504 22722
rect 7475 22717 7504 22720
rect 7551 22716 7554 22722
rect 7580 22716 7583 22742
rect 9345 22716 9348 22742
rect 9374 22736 9377 22742
rect 10251 22740 10265 22756
rect 12988 22756 13416 22770
rect 12988 22742 13002 22756
rect 10191 22737 10220 22740
rect 10191 22736 10197 22737
rect 9374 22722 10197 22736
rect 9374 22716 9377 22722
rect 10191 22720 10197 22722
rect 10214 22720 10220 22737
rect 10191 22717 10220 22720
rect 10235 22737 10265 22740
rect 10235 22720 10241 22737
rect 10258 22736 10265 22737
rect 11553 22736 11556 22742
rect 10258 22722 11556 22736
rect 10258 22720 10264 22722
rect 10235 22717 10264 22720
rect 11553 22716 11556 22722
rect 11582 22716 11585 22742
rect 12934 22737 12963 22740
rect 12934 22720 12940 22737
rect 12957 22736 12963 22737
rect 12979 22736 12982 22742
rect 12957 22722 12982 22736
rect 12957 22720 12963 22722
rect 12934 22717 12963 22720
rect 12979 22716 12982 22722
rect 13008 22716 13011 22742
rect 13026 22737 13055 22740
rect 13026 22720 13032 22737
rect 13049 22736 13055 22737
rect 13255 22736 13258 22742
rect 13049 22722 13258 22736
rect 13049 22720 13055 22722
rect 13026 22717 13055 22720
rect 13255 22716 13258 22722
rect 13284 22716 13287 22742
rect 13402 22740 13416 22756
rect 14782 22756 14980 22770
rect 15886 22756 17490 22770
rect 13394 22737 13423 22740
rect 13394 22720 13400 22737
rect 13417 22720 13423 22737
rect 13394 22717 13423 22720
rect 13624 22737 13653 22740
rect 13624 22720 13630 22737
rect 13647 22736 13653 22737
rect 13715 22736 13718 22742
rect 13647 22722 13718 22736
rect 13647 22720 13653 22722
rect 13624 22717 13653 22720
rect 13715 22716 13718 22722
rect 13744 22736 13747 22742
rect 14782 22740 14796 22756
rect 14774 22737 14803 22740
rect 13744 22722 14244 22736
rect 13744 22716 13747 22722
rect 3411 22682 3414 22708
rect 3440 22682 3443 22708
rect 7275 22682 7278 22708
rect 7304 22682 7307 22708
rect 9023 22682 9026 22708
rect 9052 22702 9055 22708
rect 9667 22702 9670 22708
rect 9052 22688 9670 22702
rect 9052 22682 9055 22688
rect 9667 22682 9670 22688
rect 9696 22702 9699 22708
rect 10036 22703 10065 22706
rect 10036 22702 10042 22703
rect 9696 22688 10042 22702
rect 9696 22682 9699 22688
rect 10036 22686 10042 22688
rect 10059 22686 10065 22703
rect 13072 22703 13101 22706
rect 13072 22702 13078 22703
rect 10036 22683 10065 22686
rect 13034 22688 13078 22702
rect 13034 22674 13048 22688
rect 13072 22686 13078 22688
rect 13095 22686 13101 22703
rect 13670 22703 13699 22706
rect 13670 22702 13676 22703
rect 13072 22683 13101 22686
rect 13632 22688 13676 22702
rect 13632 22674 13646 22688
rect 13670 22686 13676 22688
rect 13693 22686 13699 22703
rect 14230 22702 14244 22722
rect 14774 22720 14780 22737
rect 14797 22720 14803 22737
rect 14774 22717 14803 22720
rect 14819 22716 14822 22742
rect 14848 22736 14851 22742
rect 14866 22737 14895 22740
rect 14866 22736 14872 22737
rect 14848 22722 14872 22736
rect 14848 22716 14851 22722
rect 14866 22720 14872 22722
rect 14889 22720 14895 22737
rect 14866 22717 14895 22720
rect 14957 22716 14960 22742
rect 14986 22736 14989 22742
rect 15886 22740 15900 22756
rect 17487 22750 17490 22756
rect 17516 22750 17519 22776
rect 17809 22750 17812 22776
rect 17838 22770 17841 22776
rect 18324 22770 18338 22785
rect 19649 22784 19652 22790
rect 19678 22784 19681 22810
rect 17838 22756 18338 22770
rect 17838 22750 17841 22756
rect 18545 22750 18548 22776
rect 18574 22750 18577 22776
rect 21535 22750 21538 22776
rect 21564 22770 21567 22776
rect 24847 22770 24850 22776
rect 21564 22756 24850 22770
rect 21564 22750 21567 22756
rect 24847 22750 24850 22756
rect 24876 22770 24879 22776
rect 28251 22770 28254 22776
rect 24876 22756 28254 22770
rect 24876 22750 24879 22756
rect 28251 22750 28254 22756
rect 28280 22770 28283 22776
rect 28413 22771 28442 22774
rect 28413 22770 28419 22771
rect 28280 22756 28419 22770
rect 28280 22750 28283 22756
rect 28413 22754 28419 22756
rect 28436 22754 28442 22771
rect 28413 22751 28442 22754
rect 15740 22737 15769 22740
rect 15740 22736 15746 22737
rect 14986 22722 15746 22736
rect 14986 22716 14989 22722
rect 15740 22720 15746 22722
rect 15763 22720 15769 22737
rect 15740 22717 15769 22720
rect 15878 22737 15907 22740
rect 15878 22720 15884 22737
rect 15901 22720 15907 22737
rect 15878 22717 15907 22720
rect 15970 22737 15999 22740
rect 15970 22720 15976 22737
rect 15993 22736 15999 22737
rect 16245 22736 16248 22742
rect 15993 22722 16248 22736
rect 15993 22720 15999 22722
rect 15970 22717 15999 22720
rect 16245 22716 16248 22722
rect 16274 22716 16277 22742
rect 17763 22740 17766 22742
rect 17760 22717 17766 22740
rect 17763 22716 17766 22717
rect 17792 22716 17795 22742
rect 17901 22716 17904 22742
rect 17930 22736 17933 22742
rect 18554 22736 18568 22750
rect 19190 22737 19219 22740
rect 17930 22722 18154 22736
rect 18554 22722 18706 22736
rect 17930 22716 17933 22722
rect 14828 22702 14842 22716
rect 14230 22688 14842 22702
rect 13670 22683 13699 22686
rect 14911 22682 14914 22708
rect 14940 22702 14943 22708
rect 15141 22702 15144 22708
rect 14940 22688 15144 22702
rect 14940 22682 14943 22688
rect 15141 22682 15144 22688
rect 15170 22702 15173 22708
rect 16016 22703 16045 22706
rect 16016 22702 16022 22703
rect 15170 22688 16022 22702
rect 15170 22682 15173 22688
rect 16016 22686 16022 22688
rect 16039 22686 16045 22703
rect 16016 22683 16045 22686
rect 17625 22682 17628 22708
rect 17654 22682 17657 22708
rect 18140 22702 18154 22722
rect 18546 22703 18575 22706
rect 18546 22702 18552 22703
rect 18140 22688 18552 22702
rect 18546 22686 18552 22688
rect 18569 22686 18575 22703
rect 18546 22683 18575 22686
rect 18592 22703 18621 22706
rect 18637 22703 18640 22708
rect 18592 22686 18598 22703
rect 18615 22689 18640 22703
rect 18615 22686 18621 22689
rect 18592 22683 18621 22686
rect 18637 22682 18640 22689
rect 18666 22682 18669 22708
rect 18692 22706 18706 22722
rect 19190 22720 19196 22737
rect 19213 22736 19219 22737
rect 19603 22736 19606 22742
rect 19213 22722 19606 22736
rect 19213 22720 19219 22722
rect 19190 22717 19219 22720
rect 19603 22716 19606 22722
rect 19632 22716 19635 22742
rect 20064 22737 20093 22740
rect 20064 22720 20070 22737
rect 20087 22736 20093 22737
rect 21949 22736 21952 22742
rect 20087 22722 21952 22736
rect 20087 22720 20093 22722
rect 20064 22717 20093 22720
rect 21949 22716 21952 22722
rect 21978 22716 21981 22742
rect 23283 22716 23286 22742
rect 23312 22736 23315 22742
rect 23366 22737 23395 22740
rect 23366 22736 23372 22737
rect 23312 22722 23372 22736
rect 23312 22716 23315 22722
rect 23366 22720 23372 22722
rect 23389 22720 23395 22737
rect 23366 22717 23395 22720
rect 24204 22737 24233 22740
rect 24204 22720 24210 22737
rect 24227 22736 24233 22737
rect 28343 22736 28346 22742
rect 28372 22740 28375 22742
rect 28372 22737 28390 22740
rect 24227 22722 28346 22736
rect 24227 22720 24233 22722
rect 24204 22717 24233 22720
rect 18684 22703 18713 22706
rect 18684 22686 18690 22703
rect 18707 22686 18713 22703
rect 19236 22703 19265 22706
rect 19236 22702 19242 22703
rect 18684 22683 18713 22686
rect 19198 22688 19242 22702
rect 19198 22674 19212 22688
rect 19236 22686 19242 22688
rect 19259 22686 19265 22703
rect 19236 22683 19265 22686
rect 20110 22703 20139 22706
rect 20110 22686 20116 22703
rect 20133 22702 20139 22703
rect 22087 22702 22090 22708
rect 20133 22688 22090 22702
rect 20133 22686 20139 22688
rect 20110 22683 20139 22686
rect 22087 22682 22090 22688
rect 22116 22682 22119 22708
rect 23238 22703 23267 22706
rect 23238 22686 23244 22703
rect 23261 22686 23267 22703
rect 23238 22683 23267 22686
rect 13025 22648 13028 22674
rect 13054 22648 13057 22674
rect 13623 22648 13626 22674
rect 13652 22648 13655 22674
rect 19189 22648 19192 22674
rect 19218 22648 19221 22674
rect 20155 22648 20158 22674
rect 20184 22668 20187 22674
rect 20248 22669 20277 22672
rect 20248 22668 20254 22669
rect 20184 22654 20254 22668
rect 20184 22648 20187 22654
rect 20248 22652 20254 22654
rect 20271 22652 20277 22669
rect 20248 22649 20277 22652
rect 4447 22635 4476 22638
rect 4447 22618 4453 22635
rect 4470 22634 4476 22635
rect 4791 22634 4794 22640
rect 4470 22620 4794 22634
rect 4470 22618 4476 22620
rect 4447 22615 4476 22618
rect 4791 22614 4794 22620
rect 4820 22614 4823 22640
rect 8311 22635 8340 22638
rect 8311 22618 8317 22635
rect 8334 22634 8340 22635
rect 8655 22634 8658 22640
rect 8334 22620 8658 22634
rect 8334 22618 8340 22620
rect 8311 22615 8340 22618
rect 8655 22614 8658 22620
rect 8684 22614 8687 22640
rect 17717 22614 17720 22640
rect 17746 22634 17749 22640
rect 18499 22634 18502 22640
rect 17746 22620 18502 22634
rect 17746 22614 17749 22620
rect 18499 22614 18502 22620
rect 18528 22614 18531 22640
rect 18545 22614 18548 22640
rect 18574 22634 18577 22640
rect 18638 22635 18667 22638
rect 18638 22634 18644 22635
rect 18574 22620 18644 22634
rect 18574 22614 18577 22620
rect 18638 22618 18644 22620
rect 18661 22618 18667 22635
rect 23246 22634 23260 22683
rect 24157 22682 24160 22708
rect 24186 22682 24189 22708
rect 23928 22669 23957 22672
rect 23928 22652 23934 22669
rect 23951 22668 23957 22669
rect 24212 22668 24226 22717
rect 28343 22716 28346 22722
rect 28384 22720 28390 22737
rect 28372 22717 28390 22720
rect 28372 22716 28375 22717
rect 24249 22682 24252 22708
rect 24278 22702 24281 22708
rect 24296 22703 24325 22706
rect 24296 22702 24302 22703
rect 24278 22688 24302 22702
rect 24278 22682 24281 22688
rect 24296 22686 24302 22688
rect 24319 22686 24325 22703
rect 24296 22683 24325 22686
rect 28205 22682 28208 22708
rect 28234 22682 28237 22708
rect 23951 22654 24226 22668
rect 23951 22652 23957 22654
rect 23928 22649 23957 22652
rect 23329 22634 23332 22640
rect 23246 22620 23332 22634
rect 18638 22615 18667 22618
rect 23329 22614 23332 22620
rect 23358 22614 23361 22640
rect 24249 22614 24252 22640
rect 24278 22614 24281 22640
rect 29241 22635 29270 22638
rect 29241 22618 29247 22635
rect 29264 22634 29270 22635
rect 29723 22634 29726 22640
rect 29264 22620 29726 22634
rect 29264 22618 29270 22620
rect 29241 22615 29270 22618
rect 29723 22614 29726 22620
rect 29752 22614 29755 22640
rect 3036 22552 29992 22600
rect 6333 22533 6362 22536
rect 6333 22516 6339 22533
rect 6356 22532 6362 22533
rect 6401 22532 6404 22538
rect 6356 22518 6404 22532
rect 6356 22516 6362 22518
rect 6333 22513 6362 22516
rect 6401 22512 6404 22518
rect 6430 22512 6433 22538
rect 8287 22512 8290 22538
rect 8316 22532 8319 22538
rect 8702 22533 8731 22536
rect 8702 22532 8708 22533
rect 8316 22518 8708 22532
rect 8316 22512 8319 22518
rect 8702 22516 8708 22518
rect 8725 22516 8731 22533
rect 8702 22513 8731 22516
rect 17763 22512 17766 22538
rect 17792 22532 17795 22538
rect 17810 22533 17839 22536
rect 17810 22532 17816 22533
rect 17792 22518 17816 22532
rect 17792 22512 17795 22518
rect 17810 22516 17816 22518
rect 17833 22516 17839 22533
rect 17810 22513 17839 22516
rect 17901 22512 17904 22538
rect 17930 22532 17933 22538
rect 19144 22533 19173 22536
rect 19144 22532 19150 22533
rect 17930 22518 19150 22532
rect 17930 22512 17933 22518
rect 19144 22516 19150 22518
rect 19167 22516 19173 22533
rect 19144 22513 19173 22516
rect 23283 22512 23286 22538
rect 23312 22512 23315 22538
rect 4837 22498 4840 22504
rect 4739 22484 4840 22498
rect 3135 22410 3138 22436
rect 3164 22410 3167 22436
rect 3282 22431 3434 22435
rect 3282 22416 3297 22431
rect 3291 22414 3297 22416
rect 3314 22430 3434 22431
rect 3549 22430 3552 22436
rect 3314 22421 3552 22430
rect 3314 22414 3320 22421
rect 3420 22416 3552 22421
rect 3291 22411 3320 22414
rect 3549 22410 3552 22416
rect 3578 22410 3581 22436
rect 4739 22434 4753 22484
rect 4837 22478 4840 22484
rect 4866 22498 4869 22504
rect 4929 22498 4932 22504
rect 4866 22484 4932 22498
rect 4866 22478 4869 22484
rect 4929 22478 4932 22484
rect 4958 22478 4961 22504
rect 8655 22478 8658 22504
rect 8684 22498 8687 22504
rect 16429 22498 16432 22504
rect 8684 22484 8985 22498
rect 8684 22478 8687 22484
rect 4883 22464 4886 22470
rect 4875 22444 4886 22464
rect 4912 22464 4915 22470
rect 5021 22464 5024 22470
rect 4912 22450 5024 22464
rect 4912 22444 4915 22450
rect 5021 22444 5024 22450
rect 5050 22444 5053 22470
rect 7367 22444 7370 22470
rect 7396 22464 7399 22470
rect 7396 22450 7482 22464
rect 7396 22444 7399 22450
rect 4171 22431 4200 22434
rect 4171 22414 4177 22431
rect 4194 22430 4200 22431
rect 4654 22431 4683 22434
rect 4654 22430 4660 22431
rect 4194 22416 4660 22430
rect 4194 22414 4200 22416
rect 4171 22411 4200 22414
rect 4654 22414 4660 22416
rect 4677 22414 4683 22431
rect 4654 22411 4683 22414
rect 4731 22431 4760 22434
rect 4731 22414 4737 22431
rect 4754 22414 4760 22431
rect 4731 22411 4760 22414
rect 4791 22410 4794 22436
rect 4820 22434 4823 22436
rect 4820 22431 4834 22434
rect 4828 22414 4834 22431
rect 4875 22424 4889 22444
rect 4975 22434 4978 22436
rect 4966 22431 4978 22434
rect 4820 22411 4834 22414
rect 4867 22421 4896 22424
rect 4820 22410 4823 22411
rect 4867 22404 4873 22421
rect 4890 22404 4896 22421
rect 3181 22376 3184 22402
rect 3210 22396 3213 22402
rect 4867 22401 4896 22404
rect 4915 22421 4944 22424
rect 4915 22404 4921 22421
rect 4938 22419 4944 22421
rect 4938 22404 4952 22419
rect 4966 22414 4972 22431
rect 4966 22411 4978 22414
rect 4975 22410 4978 22411
rect 5004 22410 5007 22436
rect 5297 22410 5300 22436
rect 5326 22410 5329 22436
rect 5459 22431 5488 22434
rect 5459 22414 5465 22431
rect 5482 22430 5488 22431
rect 5573 22430 5576 22436
rect 5482 22416 5576 22430
rect 5482 22414 5488 22416
rect 5459 22411 5488 22414
rect 5573 22410 5576 22416
rect 5602 22410 5605 22436
rect 5619 22410 5622 22436
rect 5648 22430 5651 22436
rect 5941 22430 5944 22436
rect 5648 22416 5944 22430
rect 5648 22410 5651 22416
rect 5941 22410 5944 22416
rect 5970 22410 5973 22436
rect 7275 22410 7278 22436
rect 7304 22430 7307 22436
rect 7414 22431 7443 22434
rect 7414 22430 7420 22431
rect 7304 22416 7420 22430
rect 7304 22410 7307 22416
rect 7414 22414 7420 22416
rect 7437 22414 7443 22431
rect 7468 22430 7482 22450
rect 8333 22444 8336 22470
rect 8362 22464 8365 22470
rect 8449 22465 8478 22468
rect 8362 22450 8402 22464
rect 8362 22444 8365 22450
rect 7569 22431 7598 22434
rect 7569 22430 7575 22431
rect 7468 22416 7575 22430
rect 7414 22411 7443 22414
rect 7569 22414 7575 22416
rect 7592 22414 7598 22431
rect 8388 22430 8402 22450
rect 8449 22448 8455 22465
rect 8472 22464 8478 22465
rect 8472 22450 8770 22464
rect 8472 22448 8478 22450
rect 8449 22445 8478 22448
rect 8756 22434 8770 22450
rect 8848 22434 8875 22435
rect 8971 22434 8985 22484
rect 15863 22484 16432 22498
rect 15863 22464 15877 22484
rect 16429 22478 16432 22484
rect 16458 22478 16461 22504
rect 17625 22478 17628 22504
rect 17654 22498 17657 22504
rect 17654 22484 18384 22498
rect 17654 22478 17657 22484
rect 18370 22470 18384 22484
rect 23329 22478 23332 22504
rect 23358 22498 23361 22504
rect 23358 22484 24410 22498
rect 23358 22478 23361 22484
rect 24396 22470 24410 22484
rect 14920 22450 15877 22464
rect 8702 22431 8731 22434
rect 8702 22430 8708 22431
rect 8388 22416 8708 22430
rect 7569 22411 7598 22414
rect 8702 22414 8708 22416
rect 8725 22414 8731 22431
rect 8756 22431 8788 22434
rect 8756 22416 8765 22431
rect 8702 22411 8731 22414
rect 8759 22414 8765 22416
rect 8782 22414 8788 22431
rect 8848 22431 8882 22434
rect 8848 22430 8859 22431
rect 8759 22411 8788 22414
rect 8825 22416 8859 22430
rect 4915 22401 4952 22404
rect 3335 22397 3364 22400
rect 3335 22396 3341 22397
rect 3210 22382 3341 22396
rect 3210 22376 3213 22382
rect 3335 22380 3341 22382
rect 3358 22380 3364 22397
rect 3335 22377 3364 22380
rect 4653 22342 4656 22368
rect 4682 22342 4685 22368
rect 4745 22342 4748 22368
rect 4774 22362 4777 22368
rect 4938 22362 4952 22401
rect 5509 22397 5538 22400
rect 5509 22380 5515 22397
rect 5532 22396 5538 22397
rect 5628 22396 5642 22410
rect 5532 22382 5642 22396
rect 7422 22396 7436 22411
rect 7459 22396 7462 22402
rect 7422 22382 7462 22396
rect 5532 22380 5538 22382
rect 5509 22377 5538 22380
rect 7459 22376 7462 22382
rect 7488 22376 7491 22402
rect 7643 22400 7646 22402
rect 7625 22397 7646 22400
rect 7625 22380 7631 22397
rect 7625 22377 7646 22380
rect 7643 22376 7646 22377
rect 7672 22376 7675 22402
rect 8425 22376 8428 22402
rect 8454 22396 8457 22402
rect 8825 22396 8839 22416
rect 8853 22414 8859 22416
rect 8876 22414 8882 22431
rect 8963 22431 8992 22434
rect 8853 22411 8882 22414
rect 8915 22421 8944 22424
rect 8915 22404 8921 22421
rect 8938 22404 8944 22421
rect 8963 22414 8969 22431
rect 8986 22414 8992 22431
rect 8963 22411 8992 22414
rect 9014 22431 9043 22434
rect 9014 22414 9020 22431
rect 9037 22430 9043 22431
rect 9069 22430 9072 22436
rect 9037 22416 9072 22430
rect 9037 22414 9043 22416
rect 9014 22411 9043 22414
rect 9069 22410 9072 22416
rect 9098 22410 9101 22436
rect 13393 22410 13396 22436
rect 13422 22410 13425 22436
rect 13670 22431 13699 22434
rect 13670 22414 13676 22431
rect 13693 22430 13699 22431
rect 13715 22430 13718 22436
rect 13693 22416 13718 22430
rect 13693 22414 13699 22416
rect 13670 22411 13699 22414
rect 13715 22410 13718 22416
rect 13744 22410 13747 22436
rect 14497 22410 14500 22436
rect 14526 22430 14529 22436
rect 14920 22434 14934 22450
rect 17671 22444 17674 22470
rect 17700 22464 17703 22470
rect 17718 22465 17747 22468
rect 17718 22464 17724 22465
rect 17700 22450 17724 22464
rect 17700 22444 17703 22450
rect 17718 22448 17724 22450
rect 17741 22448 17747 22465
rect 17718 22445 17747 22448
rect 18361 22444 18364 22470
rect 18390 22464 18393 22470
rect 18454 22465 18483 22468
rect 18454 22464 18460 22465
rect 18390 22450 18460 22464
rect 18390 22444 18393 22450
rect 18454 22448 18460 22450
rect 18477 22448 18483 22465
rect 24249 22464 24252 22470
rect 18454 22445 18483 22448
rect 23292 22450 24252 22464
rect 14774 22431 14803 22434
rect 14774 22430 14780 22431
rect 14526 22416 14780 22430
rect 14526 22410 14529 22416
rect 14774 22414 14780 22416
rect 14797 22414 14803 22431
rect 14774 22411 14803 22414
rect 14912 22431 14941 22434
rect 14912 22414 14918 22431
rect 14935 22414 14941 22431
rect 14912 22411 14941 22414
rect 15049 22410 15052 22436
rect 15078 22410 15081 22436
rect 16291 22410 16294 22436
rect 16320 22410 16323 22436
rect 16430 22431 16459 22434
rect 16430 22414 16436 22431
rect 16453 22430 16459 22431
rect 16613 22430 16616 22436
rect 16453 22416 16616 22430
rect 16453 22414 16459 22416
rect 16430 22411 16459 22414
rect 16613 22410 16616 22416
rect 16642 22410 16645 22436
rect 17487 22410 17490 22436
rect 17516 22430 17519 22436
rect 17626 22431 17655 22434
rect 17626 22430 17632 22431
rect 17516 22416 17632 22430
rect 17516 22410 17519 22416
rect 17626 22414 17632 22416
rect 17649 22414 17655 22431
rect 17626 22411 17655 22414
rect 17810 22431 17839 22434
rect 17810 22414 17816 22431
rect 17833 22430 17839 22431
rect 17947 22430 17950 22436
rect 17833 22416 17950 22430
rect 17833 22414 17839 22416
rect 17810 22411 17839 22414
rect 17947 22410 17950 22416
rect 17976 22410 17979 22436
rect 21075 22410 21078 22436
rect 21104 22430 21107 22436
rect 21306 22431 21335 22434
rect 21306 22430 21312 22431
rect 21104 22416 21312 22430
rect 21104 22410 21107 22416
rect 21306 22414 21312 22416
rect 21329 22430 21335 22431
rect 21351 22430 21354 22436
rect 21329 22416 21354 22430
rect 21329 22414 21335 22416
rect 21306 22411 21335 22414
rect 21351 22410 21354 22416
rect 21380 22410 21383 22436
rect 21467 22431 21496 22434
rect 21467 22414 21473 22431
rect 21490 22430 21496 22431
rect 21627 22430 21630 22436
rect 21490 22416 21630 22430
rect 21490 22414 21496 22416
rect 21467 22411 21496 22414
rect 21627 22410 21630 22416
rect 21656 22410 21659 22436
rect 22962 22431 22991 22434
rect 22962 22414 22968 22431
rect 22985 22414 22991 22431
rect 22962 22411 22991 22414
rect 8915 22401 8944 22404
rect 8454 22382 8839 22396
rect 8454 22376 8457 22382
rect 4774 22348 4952 22362
rect 8923 22362 8937 22401
rect 18499 22376 18502 22402
rect 18528 22396 18531 22402
rect 21535 22400 21538 22402
rect 18577 22397 18606 22400
rect 18577 22396 18583 22397
rect 18528 22382 18583 22396
rect 18528 22376 18531 22382
rect 18577 22380 18583 22382
rect 18600 22380 18606 22397
rect 18577 22377 18606 22380
rect 21517 22397 21538 22400
rect 21517 22380 21523 22397
rect 21517 22377 21538 22380
rect 21535 22376 21538 22377
rect 21564 22376 21567 22402
rect 22970 22396 22984 22411
rect 23053 22410 23056 22436
rect 23082 22410 23085 22436
rect 23292 22434 23306 22450
rect 24249 22444 24252 22450
rect 24278 22444 24281 22470
rect 24387 22444 24390 22470
rect 24416 22444 24419 22470
rect 23284 22431 23313 22434
rect 23284 22414 23290 22431
rect 23307 22414 23313 22431
rect 23284 22411 23313 22414
rect 23375 22410 23378 22436
rect 23404 22410 23407 22436
rect 24525 22410 24528 22436
rect 24554 22434 24557 22436
rect 24554 22431 24572 22434
rect 24566 22414 24572 22431
rect 26963 22430 26966 22436
rect 24554 22411 24572 22414
rect 24672 22416 26966 22430
rect 24554 22410 24557 22411
rect 24341 22396 24344 22402
rect 22970 22382 24344 22396
rect 24341 22376 24344 22382
rect 24370 22376 24373 22402
rect 24433 22376 24436 22402
rect 24462 22396 24465 22402
rect 24595 22397 24624 22400
rect 24595 22396 24601 22397
rect 24462 22382 24601 22396
rect 24462 22376 24465 22382
rect 24595 22380 24601 22382
rect 24618 22396 24624 22397
rect 24672 22396 24686 22416
rect 26963 22410 26966 22416
rect 26992 22410 26995 22436
rect 24618 22382 24686 22396
rect 24618 22380 24624 22382
rect 24595 22377 24624 22380
rect 8977 22362 8980 22368
rect 8923 22348 8980 22362
rect 4774 22342 4777 22348
rect 8977 22342 8980 22348
rect 9006 22342 9009 22368
rect 13439 22342 13442 22368
rect 13468 22342 13471 22368
rect 13853 22342 13856 22368
rect 13882 22362 13885 22368
rect 13991 22362 13994 22368
rect 13882 22348 13994 22362
rect 13882 22342 13885 22348
rect 13991 22342 13994 22348
rect 14020 22362 14023 22368
rect 14820 22363 14849 22366
rect 14820 22362 14826 22363
rect 14020 22348 14826 22362
rect 14020 22342 14023 22348
rect 14820 22346 14826 22348
rect 14843 22346 14849 22363
rect 14820 22343 14849 22346
rect 15233 22342 15236 22368
rect 15262 22362 15265 22368
rect 15693 22362 15696 22368
rect 15262 22348 15696 22362
rect 15262 22342 15265 22348
rect 15693 22342 15696 22348
rect 15722 22362 15725 22368
rect 16200 22363 16229 22366
rect 16200 22362 16206 22363
rect 15722 22348 16206 22362
rect 15722 22342 15725 22348
rect 16200 22346 16206 22348
rect 16223 22346 16229 22363
rect 16200 22343 16229 22346
rect 17579 22342 17582 22368
rect 17608 22362 17611 22368
rect 17672 22363 17701 22366
rect 17672 22362 17678 22363
rect 17608 22348 17678 22362
rect 17608 22342 17611 22348
rect 17672 22346 17678 22348
rect 17695 22362 17701 22363
rect 17763 22362 17766 22368
rect 17695 22348 17766 22362
rect 17695 22346 17701 22348
rect 17672 22343 17701 22346
rect 17763 22342 17766 22348
rect 17792 22342 17795 22368
rect 22341 22363 22370 22366
rect 22341 22346 22347 22363
rect 22364 22362 22370 22363
rect 22731 22362 22734 22368
rect 22364 22348 22734 22362
rect 22364 22346 22370 22348
rect 22341 22343 22370 22346
rect 22731 22342 22734 22348
rect 22760 22342 22763 22368
rect 23007 22342 23010 22368
rect 23036 22342 23039 22368
rect 25399 22342 25402 22368
rect 25428 22366 25431 22368
rect 25428 22363 25452 22366
rect 25428 22346 25429 22363
rect 25446 22346 25452 22363
rect 25428 22343 25452 22346
rect 25428 22342 25431 22343
rect 3036 22280 29992 22328
rect 4539 22261 4568 22264
rect 4539 22244 4545 22261
rect 4562 22260 4568 22261
rect 4745 22260 4748 22266
rect 4562 22246 4748 22260
rect 4562 22244 4568 22246
rect 4539 22241 4568 22244
rect 4745 22240 4748 22246
rect 4774 22240 4777 22266
rect 8265 22261 8294 22264
rect 8265 22244 8271 22261
rect 8288 22260 8294 22261
rect 8425 22260 8428 22266
rect 8288 22246 8428 22260
rect 8288 22244 8294 22246
rect 8265 22241 8294 22244
rect 8425 22240 8428 22246
rect 8454 22240 8457 22266
rect 9621 22240 9624 22266
rect 9650 22260 9653 22266
rect 10357 22260 10360 22266
rect 9650 22246 10360 22260
rect 9650 22240 9653 22246
rect 10357 22240 10360 22246
rect 10386 22240 10389 22266
rect 14773 22240 14776 22266
rect 14802 22260 14805 22266
rect 14958 22261 14987 22264
rect 14958 22260 14964 22261
rect 14802 22246 14964 22260
rect 14802 22240 14805 22246
rect 14958 22244 14964 22246
rect 14981 22244 14987 22261
rect 14958 22241 14987 22244
rect 15141 22240 15144 22266
rect 15170 22260 15173 22266
rect 16200 22261 16229 22264
rect 16200 22260 16206 22261
rect 15170 22246 16206 22260
rect 15170 22240 15173 22246
rect 16200 22244 16206 22246
rect 16223 22244 16229 22261
rect 16200 22241 16229 22244
rect 18591 22240 18594 22266
rect 18620 22260 18623 22266
rect 23974 22261 24003 22264
rect 18620 22246 18660 22260
rect 18620 22240 18623 22246
rect 6999 22206 7002 22232
rect 7028 22226 7031 22232
rect 7437 22227 7466 22230
rect 7437 22226 7443 22227
rect 7028 22212 7443 22226
rect 7028 22206 7031 22212
rect 7437 22210 7443 22212
rect 7460 22210 7466 22227
rect 7437 22207 7466 22210
rect 9161 22206 9164 22232
rect 9190 22226 9193 22232
rect 9323 22227 9352 22230
rect 9323 22226 9329 22227
rect 9190 22212 9329 22226
rect 9190 22206 9193 22212
rect 9323 22210 9329 22212
rect 9346 22210 9352 22227
rect 16613 22226 16616 22232
rect 9323 22207 9352 22210
rect 15863 22212 16616 22226
rect 3549 22172 3552 22198
rect 3578 22192 3581 22198
rect 3659 22193 3688 22196
rect 3659 22192 3665 22193
rect 3578 22178 3665 22192
rect 3578 22172 3581 22178
rect 3659 22176 3665 22178
rect 3682 22176 3688 22193
rect 3659 22173 3688 22176
rect 3703 22193 3732 22196
rect 3703 22176 3709 22193
rect 3726 22192 3732 22193
rect 3779 22192 3782 22198
rect 3726 22178 3782 22192
rect 3726 22176 3732 22178
rect 3703 22173 3732 22176
rect 3779 22172 3782 22178
rect 3808 22192 3811 22198
rect 5205 22192 5208 22198
rect 3808 22178 5208 22192
rect 3808 22172 3811 22178
rect 5205 22172 5208 22178
rect 5234 22172 5237 22198
rect 7367 22172 7370 22198
rect 7396 22196 7399 22198
rect 7396 22193 7414 22196
rect 7408 22176 7414 22193
rect 7396 22173 7414 22176
rect 7396 22172 7399 22173
rect 9023 22172 9026 22198
rect 9052 22192 9055 22198
rect 9116 22193 9145 22196
rect 9116 22192 9122 22193
rect 9052 22178 9122 22192
rect 9052 22172 9055 22178
rect 9116 22176 9122 22178
rect 9139 22176 9145 22193
rect 9116 22173 9145 22176
rect 9277 22193 9306 22196
rect 9277 22176 9283 22193
rect 9300 22192 9306 22193
rect 9805 22192 9808 22198
rect 9300 22178 9808 22192
rect 9300 22176 9306 22178
rect 9277 22173 9306 22176
rect 9805 22172 9808 22178
rect 9834 22172 9837 22198
rect 14957 22172 14960 22198
rect 14986 22172 14989 22198
rect 15049 22172 15052 22198
rect 15078 22192 15081 22198
rect 15142 22193 15171 22196
rect 15142 22192 15148 22193
rect 15078 22178 15148 22192
rect 15078 22172 15081 22178
rect 15142 22176 15148 22178
rect 15165 22192 15171 22193
rect 15863 22192 15877 22212
rect 16613 22206 16616 22212
rect 16642 22206 16645 22232
rect 17165 22206 17168 22232
rect 17194 22226 17197 22232
rect 17533 22226 17536 22232
rect 17194 22212 17536 22226
rect 17194 22206 17197 22212
rect 17533 22206 17536 22212
rect 17562 22226 17565 22232
rect 17901 22226 17904 22232
rect 17562 22212 17904 22226
rect 17562 22206 17565 22212
rect 17901 22206 17904 22212
rect 17930 22226 17933 22232
rect 18500 22227 18529 22230
rect 17930 22212 17970 22226
rect 17930 22206 17933 22212
rect 15165 22178 15877 22192
rect 16200 22193 16229 22196
rect 15165 22176 15171 22178
rect 15142 22173 15171 22176
rect 16200 22176 16206 22193
rect 16223 22192 16229 22193
rect 16338 22193 16367 22196
rect 16223 22178 16314 22192
rect 16223 22176 16229 22178
rect 16200 22173 16229 22176
rect 3135 22138 3138 22164
rect 3164 22158 3167 22164
rect 3411 22158 3414 22164
rect 3164 22144 3414 22158
rect 3164 22138 3167 22144
rect 3411 22138 3414 22144
rect 3440 22158 3443 22164
rect 3504 22159 3533 22162
rect 3504 22158 3510 22159
rect 3440 22144 3510 22158
rect 3440 22138 3443 22144
rect 3504 22142 3510 22144
rect 3527 22142 3533 22159
rect 3504 22139 3533 22142
rect 7230 22159 7259 22162
rect 7230 22142 7236 22159
rect 7253 22142 7259 22159
rect 7230 22139 7259 22142
rect 7238 22090 7252 22139
rect 7459 22090 7462 22096
rect 7238 22076 7462 22090
rect 7459 22070 7462 22076
rect 7488 22070 7491 22096
rect 10151 22091 10180 22094
rect 10151 22074 10157 22091
rect 10174 22090 10180 22091
rect 10311 22090 10314 22096
rect 10174 22076 10314 22090
rect 10174 22074 10180 22076
rect 10151 22071 10180 22074
rect 10311 22070 10314 22076
rect 10340 22070 10343 22096
rect 16300 22090 16314 22178
rect 16338 22176 16344 22193
rect 16361 22176 16367 22193
rect 16338 22173 16367 22176
rect 17626 22193 17655 22196
rect 17626 22176 17632 22193
rect 17649 22192 17655 22193
rect 17809 22192 17812 22198
rect 17649 22178 17812 22192
rect 17649 22176 17655 22178
rect 17626 22173 17655 22176
rect 16346 22124 16360 22173
rect 17809 22172 17812 22178
rect 17838 22172 17841 22198
rect 17956 22196 17970 22212
rect 18500 22210 18506 22227
rect 18523 22226 18529 22227
rect 18545 22226 18548 22232
rect 18523 22212 18548 22226
rect 18523 22210 18529 22212
rect 18500 22207 18529 22210
rect 18545 22206 18548 22212
rect 18574 22206 18577 22232
rect 18646 22196 18660 22246
rect 23974 22244 23980 22261
rect 23997 22260 24003 22261
rect 23997 22246 26204 22260
rect 23997 22244 24003 22246
rect 23974 22241 24003 22244
rect 21305 22230 21308 22232
rect 21287 22227 21308 22230
rect 21287 22210 21293 22227
rect 21287 22207 21308 22210
rect 21305 22206 21308 22207
rect 21334 22206 21337 22232
rect 23007 22206 23010 22232
rect 23036 22226 23039 22232
rect 23407 22227 23436 22230
rect 23407 22226 23413 22227
rect 23036 22212 23413 22226
rect 23036 22206 23039 22212
rect 23407 22210 23413 22212
rect 23430 22210 23436 22227
rect 23407 22207 23436 22210
rect 17948 22193 17977 22196
rect 17948 22176 17954 22193
rect 17971 22176 17977 22193
rect 17948 22173 17977 22176
rect 18086 22193 18115 22196
rect 18086 22176 18092 22193
rect 18109 22192 18115 22193
rect 18592 22193 18621 22196
rect 18592 22192 18598 22193
rect 18109 22178 18598 22192
rect 18109 22176 18115 22178
rect 18086 22173 18115 22176
rect 18592 22176 18598 22178
rect 18615 22176 18621 22193
rect 18592 22173 18621 22176
rect 18638 22193 18667 22196
rect 18638 22176 18644 22193
rect 18661 22176 18667 22193
rect 18638 22173 18667 22176
rect 21075 22172 21078 22198
rect 21104 22172 21107 22198
rect 21237 22193 21266 22196
rect 21237 22176 21243 22193
rect 21260 22192 21266 22193
rect 21627 22192 21630 22198
rect 21260 22178 21630 22192
rect 21260 22176 21266 22178
rect 21237 22173 21266 22176
rect 21627 22172 21630 22178
rect 21656 22172 21659 22198
rect 23284 22193 23313 22196
rect 23284 22176 23290 22193
rect 23307 22192 23313 22193
rect 23329 22192 23332 22198
rect 23307 22178 23332 22192
rect 23307 22176 23313 22178
rect 23284 22173 23313 22176
rect 23329 22172 23332 22178
rect 23358 22172 23361 22198
rect 24258 22196 24272 22246
rect 24341 22206 24344 22232
rect 24370 22206 24373 22232
rect 25538 22227 25567 22230
rect 25538 22210 25544 22227
rect 25561 22226 25567 22227
rect 25629 22226 25632 22232
rect 25561 22212 25632 22226
rect 25561 22210 25567 22212
rect 25538 22207 25567 22210
rect 25629 22206 25632 22212
rect 25658 22206 25661 22232
rect 24250 22193 24279 22196
rect 24250 22176 24256 22193
rect 24273 22176 24279 22193
rect 24250 22173 24279 22176
rect 25399 22172 25402 22198
rect 25428 22172 25431 22198
rect 25492 22193 25521 22196
rect 25492 22176 25498 22193
rect 25515 22176 25521 22193
rect 25492 22173 25521 22176
rect 16384 22159 16413 22162
rect 16384 22142 16390 22159
rect 16407 22158 16413 22159
rect 16429 22158 16432 22164
rect 16407 22144 16432 22158
rect 16407 22142 16413 22144
rect 16384 22139 16413 22142
rect 16429 22138 16432 22144
rect 16458 22158 16461 22164
rect 17763 22158 17766 22164
rect 16458 22144 17766 22158
rect 16458 22138 16461 22144
rect 17763 22138 17766 22144
rect 17792 22138 17795 22164
rect 24203 22138 24206 22164
rect 24232 22138 24235 22164
rect 24295 22138 24298 22164
rect 24324 22158 24327 22164
rect 24342 22159 24371 22162
rect 24342 22158 24348 22159
rect 24324 22144 24348 22158
rect 24324 22138 24327 22144
rect 24342 22142 24348 22144
rect 24365 22142 24371 22159
rect 24342 22139 24371 22142
rect 17395 22124 17398 22130
rect 16346 22110 17398 22124
rect 17395 22104 17398 22110
rect 17424 22104 17427 22130
rect 18499 22104 18502 22130
rect 18528 22104 18531 22130
rect 25500 22124 25514 22173
rect 25583 22172 25586 22198
rect 25612 22172 25615 22198
rect 26190 22192 26204 22246
rect 26227 22206 26230 22232
rect 26256 22226 26259 22232
rect 26389 22227 26418 22230
rect 26389 22226 26395 22227
rect 26256 22212 26395 22226
rect 26256 22206 26259 22212
rect 26389 22210 26395 22212
rect 26412 22210 26418 22227
rect 26389 22207 26418 22210
rect 28463 22227 28492 22230
rect 28463 22210 28469 22227
rect 28486 22226 28492 22227
rect 28527 22226 28530 22232
rect 28486 22212 28530 22226
rect 28486 22210 28492 22212
rect 28463 22207 28492 22210
rect 28527 22206 28530 22212
rect 28556 22206 28559 22232
rect 26343 22193 26372 22196
rect 26343 22192 26349 22193
rect 26190 22178 26349 22192
rect 26343 22176 26349 22178
rect 26366 22192 26372 22193
rect 26871 22192 26874 22198
rect 26366 22178 26874 22192
rect 26366 22176 26372 22178
rect 26343 22173 26372 22176
rect 26871 22172 26874 22178
rect 26900 22172 26903 22198
rect 28205 22172 28208 22198
rect 28234 22192 28237 22198
rect 28252 22193 28281 22196
rect 28252 22192 28258 22193
rect 28234 22178 28258 22192
rect 28234 22172 28237 22178
rect 28252 22176 28258 22178
rect 28275 22176 28281 22193
rect 28252 22173 28281 22176
rect 28389 22172 28392 22198
rect 28418 22196 28421 22198
rect 28418 22193 28436 22196
rect 28430 22176 28436 22193
rect 28418 22173 28436 22176
rect 28418 22172 28421 22173
rect 26135 22138 26138 22164
rect 26164 22158 26167 22164
rect 26182 22159 26211 22162
rect 26182 22158 26188 22159
rect 26164 22144 26188 22158
rect 26164 22138 26167 22144
rect 26182 22142 26188 22144
rect 26205 22142 26211 22159
rect 26182 22139 26211 22142
rect 25500 22110 26204 22124
rect 16705 22090 16708 22096
rect 16300 22076 16708 22090
rect 16705 22070 16708 22076
rect 16734 22070 16737 22096
rect 22111 22091 22140 22094
rect 22111 22074 22117 22091
rect 22134 22090 22140 22091
rect 22639 22090 22642 22096
rect 22134 22076 22642 22090
rect 22134 22074 22140 22076
rect 22111 22071 22140 22074
rect 22639 22070 22642 22076
rect 22668 22070 22671 22096
rect 25675 22070 25678 22096
rect 25704 22070 25707 22096
rect 26190 22090 26204 22110
rect 27147 22090 27150 22096
rect 26190 22076 27150 22090
rect 27147 22070 27150 22076
rect 27176 22070 27179 22096
rect 27217 22091 27246 22094
rect 27217 22074 27223 22091
rect 27240 22090 27246 22091
rect 28021 22090 28024 22096
rect 27240 22076 28024 22090
rect 27240 22074 27246 22076
rect 27217 22071 27246 22074
rect 28021 22070 28024 22076
rect 28050 22070 28053 22096
rect 29287 22091 29316 22094
rect 29287 22074 29293 22091
rect 29310 22090 29316 22091
rect 29539 22090 29542 22096
rect 29310 22076 29542 22090
rect 29310 22074 29316 22076
rect 29287 22071 29316 22074
rect 29539 22070 29542 22076
rect 29568 22070 29571 22096
rect 3036 22008 29992 22056
rect 5297 21988 5300 21994
rect 5168 21974 5300 21988
rect 4929 21866 4932 21892
rect 4958 21886 4961 21892
rect 5168 21890 5182 21974
rect 5297 21968 5300 21974
rect 5326 21968 5329 21994
rect 5343 21968 5346 21994
rect 5372 21988 5375 21994
rect 5711 21988 5714 21994
rect 5372 21974 5714 21988
rect 5372 21968 5375 21974
rect 5711 21968 5714 21974
rect 5740 21988 5743 21994
rect 9713 21988 9716 21994
rect 5740 21974 9716 21988
rect 5740 21968 5743 21974
rect 9713 21968 9716 21974
rect 9742 21968 9745 21994
rect 15863 21974 17096 21988
rect 6195 21921 6224 21924
rect 6195 21904 6201 21921
rect 6218 21920 6224 21921
rect 6631 21920 6634 21926
rect 6218 21906 6516 21920
rect 6218 21904 6224 21906
rect 6195 21901 6224 21904
rect 5160 21887 5189 21890
rect 5160 21886 5166 21887
rect 4958 21872 5166 21886
rect 4958 21866 4961 21872
rect 5160 21870 5166 21872
rect 5183 21870 5189 21887
rect 5160 21867 5189 21870
rect 5321 21887 5350 21890
rect 5321 21870 5327 21887
rect 5344 21886 5350 21887
rect 5481 21886 5484 21892
rect 5344 21872 5484 21886
rect 5344 21870 5350 21872
rect 5321 21867 5350 21870
rect 5481 21866 5484 21872
rect 5510 21866 5513 21892
rect 6447 21866 6450 21892
rect 6476 21866 6479 21892
rect 6502 21890 6516 21906
rect 6594 21906 6634 21920
rect 6594 21890 6608 21906
rect 6631 21900 6634 21906
rect 6660 21900 6663 21926
rect 6494 21887 6523 21890
rect 6494 21870 6500 21887
rect 6517 21870 6523 21887
rect 6494 21867 6523 21870
rect 6586 21887 6615 21890
rect 6586 21870 6592 21887
rect 6609 21870 6615 21887
rect 6586 21867 6615 21870
rect 6678 21887 6707 21890
rect 6678 21870 6684 21887
rect 6701 21886 6707 21887
rect 6723 21886 6726 21892
rect 6701 21872 6726 21886
rect 6701 21870 6707 21872
rect 6678 21867 6707 21870
rect 6723 21866 6726 21872
rect 6752 21866 6755 21892
rect 10173 21866 10176 21892
rect 10202 21866 10205 21892
rect 10265 21866 10268 21892
rect 10294 21866 10297 21892
rect 10311 21866 10314 21892
rect 10340 21866 10343 21892
rect 10357 21866 10360 21892
rect 10386 21866 10389 21892
rect 11324 21887 11353 21890
rect 11324 21870 11330 21887
rect 11347 21886 11353 21887
rect 11369 21886 11372 21892
rect 11347 21872 11372 21886
rect 11347 21870 11353 21872
rect 11324 21867 11353 21870
rect 11369 21866 11372 21872
rect 11398 21866 11401 21892
rect 11461 21866 11464 21892
rect 11490 21890 11493 21892
rect 11490 21887 11508 21890
rect 11502 21870 11508 21887
rect 11490 21867 11508 21870
rect 14406 21887 14435 21890
rect 14406 21870 14412 21887
rect 14429 21886 14435 21887
rect 14497 21886 14500 21892
rect 14429 21872 14500 21886
rect 14429 21870 14435 21872
rect 14406 21867 14435 21870
rect 11490 21866 11493 21867
rect 14497 21866 14500 21872
rect 14526 21866 14529 21892
rect 14544 21887 14573 21890
rect 14544 21870 14550 21887
rect 14567 21870 14573 21887
rect 14544 21867 14573 21870
rect 5205 21832 5208 21858
rect 5234 21852 5237 21858
rect 5367 21853 5396 21856
rect 5367 21852 5373 21853
rect 5234 21838 5373 21852
rect 5234 21832 5237 21838
rect 5367 21836 5373 21838
rect 5390 21836 5396 21853
rect 5367 21833 5396 21836
rect 6631 21832 6634 21858
rect 6660 21832 6663 21858
rect 11553 21856 11556 21858
rect 11535 21853 11556 21856
rect 11535 21836 11541 21853
rect 11535 21833 11556 21836
rect 11553 21832 11556 21833
rect 11582 21832 11585 21858
rect 14552 21852 14566 21867
rect 14957 21866 14960 21892
rect 14986 21866 14989 21892
rect 15142 21887 15171 21890
rect 15142 21870 15148 21887
rect 15165 21886 15171 21887
rect 15863 21886 15877 21974
rect 16484 21940 17050 21954
rect 16484 21890 16498 21940
rect 15165 21872 15877 21886
rect 16338 21887 16367 21890
rect 15165 21870 15171 21872
rect 15142 21867 15171 21870
rect 16338 21870 16344 21887
rect 16361 21870 16367 21887
rect 16338 21867 16367 21870
rect 16476 21887 16505 21890
rect 16476 21870 16482 21887
rect 16499 21870 16505 21887
rect 16476 21867 16505 21870
rect 16522 21887 16551 21890
rect 16522 21870 16528 21887
rect 16545 21886 16551 21887
rect 16613 21886 16616 21892
rect 16545 21872 16616 21886
rect 16545 21870 16551 21872
rect 16522 21867 16551 21870
rect 15150 21852 15164 21867
rect 14552 21838 15164 21852
rect 16346 21852 16360 21867
rect 16613 21866 16616 21872
rect 16642 21866 16645 21892
rect 17036 21890 17050 21940
rect 17082 21924 17096 21974
rect 17487 21968 17490 21994
rect 17516 21988 17519 21994
rect 17672 21989 17701 21992
rect 17672 21988 17678 21989
rect 17516 21974 17678 21988
rect 17516 21968 17519 21974
rect 17672 21972 17678 21974
rect 17695 21972 17701 21989
rect 17672 21969 17701 21972
rect 23053 21968 23056 21994
rect 23082 21988 23085 21994
rect 23238 21989 23267 21992
rect 23238 21988 23244 21989
rect 23082 21974 23244 21988
rect 23082 21968 23085 21974
rect 23238 21972 23244 21974
rect 23261 21972 23267 21989
rect 25583 21988 25586 21994
rect 23238 21969 23267 21972
rect 23292 21974 25586 21988
rect 17074 21921 17103 21924
rect 17074 21904 17080 21921
rect 17097 21920 17103 21921
rect 17717 21920 17720 21926
rect 17097 21906 17720 21920
rect 17097 21904 17103 21906
rect 17074 21901 17103 21904
rect 17717 21900 17720 21906
rect 17746 21900 17749 21926
rect 17901 21900 17904 21926
rect 17930 21900 17933 21926
rect 19373 21900 19376 21926
rect 19402 21920 19405 21926
rect 19512 21921 19541 21924
rect 19512 21920 19518 21921
rect 19402 21906 19518 21920
rect 19402 21900 19405 21906
rect 19512 21904 19518 21906
rect 19535 21904 19541 21921
rect 19512 21901 19541 21904
rect 21075 21900 21078 21926
rect 21104 21920 21107 21926
rect 21214 21921 21243 21924
rect 21214 21920 21220 21921
rect 21104 21906 21220 21920
rect 21104 21900 21107 21906
rect 21214 21904 21220 21906
rect 21237 21904 21243 21921
rect 21214 21901 21243 21904
rect 22249 21921 22278 21924
rect 22249 21904 22255 21921
rect 22272 21920 22278 21921
rect 22272 21906 22570 21920
rect 22272 21904 22278 21906
rect 22249 21901 22278 21904
rect 16890 21887 16919 21890
rect 16890 21870 16896 21887
rect 16913 21870 16919 21887
rect 16890 21867 16919 21870
rect 17028 21887 17057 21890
rect 17028 21870 17034 21887
rect 17051 21886 17057 21887
rect 17533 21886 17536 21892
rect 17051 21872 17536 21886
rect 17051 21870 17057 21872
rect 17028 21867 17057 21870
rect 16898 21852 16912 21867
rect 17533 21866 17536 21872
rect 17562 21866 17565 21892
rect 17809 21866 17812 21892
rect 17838 21886 17841 21892
rect 17856 21887 17885 21890
rect 17856 21886 17862 21887
rect 17838 21872 17862 21886
rect 17838 21866 17841 21872
rect 17856 21870 17862 21872
rect 17879 21870 17885 21887
rect 17856 21867 17885 21870
rect 19673 21887 19702 21890
rect 19673 21870 19679 21887
rect 19696 21886 19702 21887
rect 19787 21886 19790 21892
rect 19696 21872 19790 21886
rect 19696 21870 19702 21872
rect 19673 21867 19702 21870
rect 19787 21866 19790 21872
rect 19816 21866 19819 21892
rect 21121 21886 21124 21892
rect 19842 21872 21124 21886
rect 17818 21852 17832 21866
rect 16346 21838 17832 21852
rect 19723 21853 19752 21856
rect 19723 21836 19729 21853
rect 19746 21852 19752 21853
rect 19842 21852 19856 21872
rect 21121 21866 21124 21872
rect 21150 21866 21153 21892
rect 21375 21887 21404 21890
rect 21375 21870 21381 21887
rect 21398 21886 21404 21887
rect 21627 21886 21630 21892
rect 21398 21872 21630 21886
rect 21398 21870 21404 21872
rect 21375 21867 21404 21870
rect 21627 21866 21630 21872
rect 21656 21866 21659 21892
rect 22501 21866 22504 21892
rect 22530 21866 22533 21892
rect 22556 21890 22570 21906
rect 22731 21900 22734 21926
rect 22760 21920 22763 21926
rect 23292 21920 23306 21974
rect 25583 21968 25586 21974
rect 25612 21988 25615 21994
rect 26181 21988 26184 21994
rect 25612 21974 26184 21988
rect 25612 21968 25615 21974
rect 26181 21968 26184 21974
rect 26210 21968 26213 21994
rect 27377 21968 27380 21994
rect 27406 21988 27409 21994
rect 28022 21989 28051 21992
rect 28022 21988 28028 21989
rect 27406 21974 28028 21988
rect 27406 21968 27409 21974
rect 28022 21972 28028 21974
rect 28045 21972 28051 21989
rect 28022 21969 28051 21972
rect 25629 21934 25632 21960
rect 25658 21954 25661 21960
rect 25722 21955 25751 21958
rect 25722 21954 25728 21955
rect 25658 21940 25728 21954
rect 25658 21934 25661 21940
rect 25722 21938 25728 21940
rect 25745 21938 25751 21955
rect 25722 21935 25751 21938
rect 27769 21955 27798 21958
rect 27769 21938 27775 21955
rect 27792 21954 27798 21955
rect 27792 21940 28296 21954
rect 27792 21938 27798 21940
rect 27769 21935 27798 21938
rect 22760 21900 22767 21920
rect 22556 21887 22588 21890
rect 22556 21872 22565 21887
rect 22559 21870 22565 21872
rect 22582 21870 22588 21887
rect 22559 21867 22588 21870
rect 22639 21866 22642 21892
rect 22668 21890 22671 21892
rect 22668 21887 22682 21890
rect 22676 21870 22682 21887
rect 22753 21880 22767 21900
rect 23200 21906 23306 21920
rect 22814 21887 22843 21890
rect 22668 21867 22682 21870
rect 22701 21877 22730 21880
rect 22668 21866 22671 21867
rect 22701 21860 22707 21877
rect 22724 21860 22730 21877
rect 21443 21856 21446 21858
rect 19746 21838 19856 21852
rect 21425 21853 21446 21856
rect 19746 21836 19752 21838
rect 19723 21833 19752 21836
rect 21425 21836 21431 21853
rect 21425 21833 21446 21836
rect 21443 21832 21446 21833
rect 21472 21832 21475 21858
rect 22317 21832 22320 21858
rect 22346 21852 22349 21858
rect 22701 21857 22730 21860
rect 22749 21877 22778 21880
rect 22749 21860 22755 21877
rect 22772 21860 22778 21877
rect 22814 21870 22820 21887
rect 22837 21886 22843 21887
rect 23007 21886 23010 21892
rect 22837 21872 23010 21886
rect 22837 21870 22843 21872
rect 22814 21867 22843 21870
rect 23007 21866 23010 21872
rect 23036 21886 23039 21892
rect 23200 21886 23214 21906
rect 24387 21900 24390 21926
rect 24416 21920 24419 21926
rect 24434 21921 24463 21924
rect 24434 21920 24440 21921
rect 24416 21906 24440 21920
rect 24416 21900 24419 21906
rect 24434 21904 24440 21906
rect 24457 21904 24463 21921
rect 26227 21920 26230 21926
rect 24434 21901 24463 21904
rect 25523 21906 26230 21920
rect 23036 21872 23214 21886
rect 23036 21866 23039 21872
rect 23237 21866 23240 21892
rect 23266 21866 23269 21892
rect 23329 21886 23332 21892
rect 23292 21872 23332 21886
rect 22749 21857 22778 21860
rect 22346 21838 22570 21852
rect 22346 21832 22349 21838
rect 6539 21798 6542 21824
rect 6568 21798 6571 21824
rect 10450 21819 10479 21822
rect 10450 21802 10456 21819
rect 10473 21818 10479 21819
rect 10587 21818 10590 21824
rect 10473 21804 10590 21818
rect 10473 21802 10479 21804
rect 10450 21799 10479 21802
rect 10587 21798 10590 21804
rect 10616 21798 10619 21824
rect 12359 21819 12388 21822
rect 12359 21802 12365 21819
rect 12382 21818 12388 21819
rect 12427 21818 12430 21824
rect 12382 21804 12430 21818
rect 12382 21802 12388 21804
rect 12359 21799 12388 21802
rect 12427 21798 12430 21804
rect 12456 21798 12459 21824
rect 14083 21798 14086 21824
rect 14112 21818 14115 21824
rect 14314 21819 14343 21822
rect 14314 21818 14320 21819
rect 14112 21804 14320 21818
rect 14112 21798 14115 21804
rect 14314 21802 14320 21804
rect 14337 21802 14343 21819
rect 14314 21799 14343 21802
rect 14359 21798 14362 21824
rect 14388 21818 14391 21824
rect 14912 21819 14941 21822
rect 14912 21818 14918 21819
rect 14388 21804 14918 21818
rect 14388 21798 14391 21804
rect 14912 21802 14918 21804
rect 14935 21802 14941 21819
rect 14912 21799 14941 21802
rect 16337 21798 16340 21824
rect 16366 21798 16369 21824
rect 16429 21798 16432 21824
rect 16458 21818 16461 21824
rect 16521 21818 16524 21824
rect 16458 21804 16524 21818
rect 16458 21798 16461 21804
rect 16521 21798 16524 21804
rect 16550 21818 16553 21824
rect 16890 21819 16919 21822
rect 16890 21818 16896 21819
rect 16550 21804 16896 21818
rect 16550 21798 16553 21804
rect 16890 21802 16896 21804
rect 16913 21802 16919 21819
rect 16890 21799 16919 21802
rect 20547 21819 20576 21822
rect 20547 21802 20553 21819
rect 20570 21818 20576 21819
rect 20661 21818 20664 21824
rect 20570 21804 20664 21818
rect 20570 21802 20576 21804
rect 20547 21799 20576 21802
rect 20661 21798 20664 21804
rect 20690 21798 20693 21824
rect 22501 21798 22504 21824
rect 22530 21798 22533 21824
rect 22556 21818 22570 21838
rect 22709 21818 22723 21857
rect 23191 21832 23194 21858
rect 23220 21852 23223 21858
rect 23292 21852 23306 21872
rect 23329 21866 23332 21872
rect 23358 21866 23361 21892
rect 25523 21886 25537 21906
rect 26227 21900 26230 21906
rect 26256 21900 26259 21926
rect 28282 21896 28296 21940
rect 28275 21893 28304 21896
rect 24672 21872 25537 21886
rect 24672 21858 24686 21872
rect 25675 21866 25678 21892
rect 25704 21886 25707 21892
rect 25722 21887 25751 21890
rect 25722 21886 25728 21887
rect 25704 21872 25728 21886
rect 25704 21866 25707 21872
rect 25722 21870 25728 21872
rect 25745 21870 25751 21887
rect 25722 21867 25751 21870
rect 25859 21866 25862 21892
rect 25888 21866 25891 21892
rect 26135 21866 26138 21892
rect 26164 21886 26167 21892
rect 26734 21887 26763 21890
rect 26734 21886 26740 21887
rect 26164 21872 26740 21886
rect 26164 21866 26167 21872
rect 26734 21870 26740 21872
rect 26757 21870 26763 21887
rect 26734 21867 26763 21870
rect 26871 21866 26874 21892
rect 26900 21890 26903 21892
rect 26900 21887 26918 21890
rect 26912 21870 26918 21887
rect 26900 21867 26918 21870
rect 26900 21866 26903 21867
rect 28021 21866 28024 21892
rect 28050 21866 28053 21892
rect 28067 21866 28070 21892
rect 28096 21890 28099 21892
rect 28096 21887 28108 21890
rect 28102 21870 28108 21887
rect 28096 21867 28108 21870
rect 28096 21866 28099 21867
rect 28159 21866 28162 21892
rect 28188 21890 28191 21892
rect 28188 21887 28209 21890
rect 28203 21870 28209 21887
rect 28188 21867 28209 21870
rect 28228 21877 28257 21880
rect 28188 21866 28191 21867
rect 28228 21860 28234 21877
rect 28251 21860 28257 21877
rect 28275 21876 28281 21893
rect 28298 21876 28304 21893
rect 28343 21890 28346 21892
rect 28275 21873 28304 21876
rect 28334 21887 28346 21890
rect 28334 21870 28340 21887
rect 28334 21867 28346 21870
rect 28343 21866 28346 21867
rect 28372 21866 28375 21892
rect 23220 21838 23306 21852
rect 23220 21832 23223 21838
rect 24479 21832 24482 21858
rect 24508 21852 24511 21858
rect 24663 21856 24666 21858
rect 24594 21853 24623 21856
rect 24594 21852 24600 21853
rect 24508 21838 24600 21852
rect 24508 21832 24511 21838
rect 24594 21836 24600 21838
rect 24617 21836 24623 21853
rect 24594 21833 24623 21836
rect 24645 21853 24666 21856
rect 24645 21836 24651 21853
rect 24645 21833 24666 21836
rect 24663 21832 24666 21833
rect 24692 21832 24695 21858
rect 26963 21856 26966 21858
rect 26945 21853 26966 21856
rect 26945 21836 26951 21853
rect 26945 21833 26966 21836
rect 26963 21832 26966 21833
rect 26992 21832 26995 21858
rect 28228 21857 28257 21860
rect 22556 21804 22723 21818
rect 25469 21819 25498 21822
rect 25469 21802 25475 21819
rect 25492 21818 25498 21819
rect 25814 21819 25843 21822
rect 25814 21818 25820 21819
rect 25492 21804 25820 21818
rect 25492 21802 25498 21804
rect 25469 21799 25498 21802
rect 25814 21802 25820 21804
rect 25837 21802 25843 21819
rect 25814 21799 25843 21802
rect 27193 21798 27196 21824
rect 27222 21818 27225 21824
rect 28229 21818 28243 21857
rect 27222 21804 28243 21818
rect 27222 21798 27225 21804
rect 3036 21736 29992 21784
rect 4792 21717 4821 21720
rect 4792 21700 4798 21717
rect 4815 21716 4821 21717
rect 6447 21716 6450 21722
rect 4815 21702 6450 21716
rect 4815 21700 4821 21702
rect 4792 21697 4821 21700
rect 6447 21696 6450 21702
rect 6476 21696 6479 21722
rect 15509 21696 15512 21722
rect 15538 21716 15541 21722
rect 15538 21702 16038 21716
rect 15538 21696 15541 21702
rect 3457 21662 3460 21688
rect 3486 21682 3489 21688
rect 3641 21686 3644 21688
rect 3623 21683 3644 21686
rect 3623 21682 3629 21683
rect 3486 21668 3629 21682
rect 3486 21662 3489 21668
rect 3623 21666 3629 21668
rect 3623 21663 3644 21666
rect 3641 21662 3644 21663
rect 3670 21662 3673 21688
rect 4653 21662 4656 21688
rect 4682 21682 4685 21688
rect 4746 21683 4775 21686
rect 4746 21682 4752 21683
rect 4682 21668 4752 21682
rect 4682 21662 4685 21668
rect 4746 21666 4752 21668
rect 4769 21666 4775 21683
rect 4746 21663 4775 21666
rect 7229 21662 7232 21688
rect 7258 21682 7261 21688
rect 7436 21683 7465 21686
rect 7436 21682 7442 21683
rect 7258 21668 7442 21682
rect 7258 21662 7261 21668
rect 7436 21666 7442 21668
rect 7459 21666 7465 21683
rect 7436 21663 7465 21666
rect 7487 21683 7516 21686
rect 7487 21666 7493 21683
rect 7510 21682 7516 21683
rect 7510 21668 7620 21682
rect 7510 21666 7516 21668
rect 7487 21663 7516 21666
rect 7606 21654 7620 21668
rect 8517 21662 8520 21688
rect 8546 21682 8549 21688
rect 9897 21686 9900 21688
rect 9879 21683 9900 21686
rect 9879 21682 9885 21683
rect 8546 21668 9885 21682
rect 8546 21662 8549 21668
rect 9879 21666 9885 21668
rect 9879 21663 9900 21666
rect 9897 21662 9900 21663
rect 9926 21662 9929 21688
rect 11875 21686 11878 21688
rect 11857 21683 11878 21686
rect 11857 21666 11863 21683
rect 11857 21663 11878 21666
rect 11875 21662 11878 21663
rect 11904 21662 11907 21688
rect 12657 21662 12660 21688
rect 12686 21682 12689 21688
rect 14543 21686 14546 21688
rect 13302 21683 13331 21686
rect 13302 21682 13308 21683
rect 12686 21668 13308 21682
rect 12686 21662 12689 21668
rect 13302 21666 13308 21668
rect 13325 21666 13331 21683
rect 13302 21663 13331 21666
rect 14525 21683 14546 21686
rect 14525 21666 14531 21683
rect 14525 21663 14546 21666
rect 14543 21662 14546 21663
rect 14572 21662 14575 21688
rect 3549 21628 3552 21654
rect 3578 21652 3581 21654
rect 3578 21649 3596 21652
rect 3590 21632 3596 21649
rect 3578 21629 3596 21632
rect 3578 21628 3581 21629
rect 4837 21628 4840 21654
rect 4866 21628 4869 21654
rect 4883 21628 4886 21654
rect 4912 21628 4915 21654
rect 6402 21649 6431 21652
rect 6402 21632 6408 21649
rect 6425 21632 6431 21649
rect 6402 21629 6431 21632
rect 3411 21594 3414 21620
rect 3440 21594 3443 21620
rect 6410 21614 6424 21629
rect 6493 21628 6496 21654
rect 6522 21628 6525 21654
rect 6539 21628 6542 21654
rect 6568 21648 6571 21654
rect 6632 21649 6661 21652
rect 6632 21648 6638 21649
rect 6568 21634 6638 21648
rect 6568 21628 6571 21634
rect 6632 21632 6638 21634
rect 6655 21632 6661 21649
rect 6632 21629 6661 21632
rect 7597 21628 7600 21654
rect 7626 21628 7629 21654
rect 9667 21628 9670 21654
rect 9696 21628 9699 21654
rect 9805 21628 9808 21654
rect 9834 21652 9837 21654
rect 9834 21649 9852 21652
rect 9846 21632 9852 21649
rect 9834 21629 9852 21632
rect 9834 21628 9837 21629
rect 11461 21628 11464 21654
rect 11490 21648 11493 21654
rect 11801 21649 11830 21652
rect 11801 21648 11807 21649
rect 11490 21634 11807 21648
rect 11490 21628 11493 21634
rect 11801 21632 11807 21634
rect 11824 21632 11830 21649
rect 11801 21629 11830 21632
rect 12703 21628 12706 21654
rect 12732 21648 12735 21654
rect 13026 21649 13055 21652
rect 13026 21648 13032 21649
rect 12732 21634 13032 21648
rect 12732 21628 12735 21634
rect 13026 21632 13032 21634
rect 13049 21632 13055 21649
rect 13026 21629 13055 21632
rect 13071 21628 13074 21654
rect 13100 21628 13103 21654
rect 14221 21628 14224 21654
rect 14250 21648 14253 21654
rect 14469 21649 14498 21652
rect 14469 21648 14475 21649
rect 14250 21634 14475 21648
rect 14250 21628 14253 21634
rect 14469 21632 14475 21634
rect 14492 21632 14498 21649
rect 14469 21629 14498 21632
rect 15831 21628 15834 21654
rect 15860 21628 15863 21654
rect 16024 21652 16038 21702
rect 18223 21696 18226 21722
rect 18252 21696 18255 21722
rect 21443 21696 21446 21722
rect 21472 21716 21475 21722
rect 21673 21716 21676 21722
rect 21472 21702 21676 21716
rect 21472 21696 21475 21702
rect 21673 21696 21676 21702
rect 21702 21696 21705 21722
rect 22455 21696 22458 21722
rect 22484 21716 22487 21722
rect 22547 21716 22550 21722
rect 22484 21702 22550 21716
rect 22484 21696 22487 21702
rect 22547 21696 22550 21702
rect 22576 21716 22579 21722
rect 25859 21716 25862 21722
rect 22576 21702 25862 21716
rect 22576 21696 22579 21702
rect 25859 21696 25862 21702
rect 25888 21696 25891 21722
rect 27171 21717 27200 21720
rect 27171 21700 27177 21717
rect 27194 21716 27200 21717
rect 28159 21716 28162 21722
rect 27194 21702 28162 21716
rect 27194 21700 27200 21702
rect 27171 21697 27200 21700
rect 28159 21696 28162 21702
rect 28188 21696 28191 21722
rect 16705 21662 16708 21688
rect 16734 21682 16737 21688
rect 16734 21668 17556 21682
rect 16734 21662 16737 21668
rect 15878 21649 15907 21652
rect 15878 21632 15884 21649
rect 15901 21632 15907 21649
rect 15878 21629 15907 21632
rect 16016 21649 16045 21652
rect 16016 21632 16022 21649
rect 16039 21632 16045 21649
rect 16016 21629 16045 21632
rect 6410 21600 6516 21614
rect 4699 21560 4702 21586
rect 4728 21580 4731 21586
rect 4728 21566 6217 21580
rect 4728 21560 4731 21566
rect 4447 21547 4476 21550
rect 4447 21530 4453 21547
rect 4470 21546 4476 21547
rect 4791 21546 4794 21552
rect 4470 21532 4794 21546
rect 4470 21530 4476 21532
rect 4447 21527 4476 21530
rect 4791 21526 4794 21532
rect 4820 21526 4823 21552
rect 6203 21546 6217 21566
rect 6448 21547 6477 21550
rect 6448 21546 6454 21547
rect 6203 21532 6454 21546
rect 6448 21530 6454 21532
rect 6471 21530 6477 21547
rect 6502 21546 6516 21600
rect 7275 21594 7278 21620
rect 7304 21594 7307 21620
rect 11415 21594 11418 21620
rect 11444 21614 11447 21620
rect 11646 21615 11675 21618
rect 11646 21614 11652 21615
rect 11444 21600 11652 21614
rect 11444 21594 11447 21600
rect 11646 21598 11652 21600
rect 11669 21598 11675 21615
rect 11646 21595 11675 21598
rect 14175 21594 14178 21620
rect 14204 21614 14207 21620
rect 14314 21615 14343 21618
rect 14314 21614 14320 21615
rect 14204 21600 14320 21614
rect 14204 21594 14207 21600
rect 14314 21598 14320 21600
rect 14337 21598 14343 21615
rect 14314 21595 14343 21598
rect 15349 21615 15378 21618
rect 15349 21598 15355 21615
rect 15372 21614 15378 21615
rect 15886 21614 15900 21629
rect 16153 21628 16156 21654
rect 16182 21628 16185 21654
rect 16245 21628 16248 21654
rect 16274 21628 16277 21654
rect 17395 21628 17398 21654
rect 17424 21648 17427 21654
rect 17488 21649 17517 21652
rect 17488 21648 17494 21649
rect 17424 21634 17494 21648
rect 17424 21628 17427 21634
rect 17488 21632 17494 21634
rect 17511 21632 17517 21649
rect 17542 21648 17556 21668
rect 17717 21662 17720 21688
rect 17746 21662 17749 21688
rect 21682 21682 21696 21696
rect 24663 21682 24666 21688
rect 17864 21668 18338 21682
rect 21682 21668 24666 21682
rect 17810 21649 17839 21652
rect 17810 21648 17816 21649
rect 17542 21634 17816 21648
rect 17488 21629 17517 21632
rect 17810 21632 17816 21634
rect 17833 21632 17839 21649
rect 17810 21629 17839 21632
rect 15372 21600 15900 21614
rect 16162 21614 16176 21628
rect 16429 21614 16432 21620
rect 16162 21600 16432 21614
rect 15372 21598 15378 21600
rect 15349 21595 15378 21598
rect 16429 21594 16432 21600
rect 16458 21594 16461 21620
rect 17496 21614 17510 21629
rect 17864 21614 17878 21668
rect 18324 21652 18338 21668
rect 24663 21662 24666 21668
rect 24692 21662 24695 21688
rect 26365 21686 26368 21688
rect 26347 21683 26368 21686
rect 26347 21666 26353 21683
rect 26347 21663 26368 21666
rect 26365 21662 26368 21663
rect 26394 21662 26397 21688
rect 28435 21686 28438 21688
rect 28417 21683 28438 21686
rect 28417 21666 28423 21683
rect 28417 21663 28438 21666
rect 28435 21662 28438 21663
rect 28464 21662 28467 21688
rect 29241 21683 29270 21686
rect 29241 21666 29247 21683
rect 29264 21682 29270 21683
rect 29264 21668 29637 21682
rect 29264 21666 29270 21668
rect 29241 21663 29270 21666
rect 17948 21649 17977 21652
rect 17948 21632 17954 21649
rect 17971 21648 17977 21649
rect 18178 21649 18207 21652
rect 18178 21648 18184 21649
rect 17971 21634 18184 21648
rect 17971 21632 17977 21634
rect 17948 21629 17977 21632
rect 18178 21632 18184 21634
rect 18201 21632 18207 21649
rect 18178 21629 18207 21632
rect 18316 21649 18345 21652
rect 18316 21632 18322 21649
rect 18339 21632 18345 21649
rect 18316 21629 18345 21632
rect 26297 21649 26326 21652
rect 26297 21632 26303 21649
rect 26320 21648 26326 21649
rect 26871 21648 26874 21654
rect 26320 21634 26874 21648
rect 26320 21632 26326 21634
rect 26297 21629 26326 21632
rect 26871 21628 26874 21634
rect 26900 21628 26903 21654
rect 28205 21628 28208 21654
rect 28234 21628 28237 21654
rect 28343 21628 28346 21654
rect 28372 21652 28375 21654
rect 28372 21649 28390 21652
rect 28384 21632 28390 21649
rect 28372 21629 28390 21632
rect 28372 21628 28375 21629
rect 29355 21628 29358 21654
rect 29384 21648 29387 21654
rect 29494 21649 29523 21652
rect 29494 21648 29500 21649
rect 29384 21634 29500 21648
rect 29384 21628 29387 21634
rect 29494 21632 29500 21634
rect 29517 21632 29523 21649
rect 29494 21629 29523 21632
rect 29539 21628 29542 21654
rect 29568 21652 29571 21654
rect 29568 21649 29580 21652
rect 29574 21632 29580 21649
rect 29623 21648 29637 21668
rect 29723 21662 29726 21688
rect 29752 21682 29755 21688
rect 29752 21668 29792 21682
rect 29752 21662 29755 21668
rect 29652 21649 29681 21652
rect 29652 21648 29658 21649
rect 29623 21634 29658 21648
rect 29568 21629 29580 21632
rect 29652 21632 29658 21634
rect 29675 21632 29681 21649
rect 29778 21647 29792 21668
rect 29815 21652 29818 21654
rect 29652 21629 29681 21632
rect 29707 21644 29736 21647
rect 29568 21628 29571 21629
rect 29707 21627 29713 21644
rect 29730 21627 29736 21644
rect 29707 21624 29736 21627
rect 29755 21644 29792 21647
rect 29755 21627 29761 21644
rect 29778 21628 29792 21644
rect 29806 21649 29818 21652
rect 29806 21632 29812 21649
rect 29806 21629 29818 21632
rect 29815 21628 29818 21629
rect 29844 21628 29847 21654
rect 29778 21627 29784 21628
rect 29755 21624 29784 21627
rect 17496 21600 17878 21614
rect 17901 21594 17904 21620
rect 17930 21614 17933 21620
rect 18408 21615 18437 21618
rect 18408 21614 18414 21615
rect 17930 21600 18414 21614
rect 17930 21594 17933 21600
rect 18408 21598 18414 21600
rect 18431 21598 18437 21615
rect 18408 21595 18437 21598
rect 25537 21594 25540 21620
rect 25566 21614 25569 21620
rect 26135 21614 26138 21620
rect 25566 21600 26138 21614
rect 25566 21594 25569 21600
rect 26135 21594 26138 21600
rect 26164 21594 26167 21620
rect 12934 21581 12963 21584
rect 12934 21580 12940 21581
rect 12482 21566 12940 21580
rect 7643 21546 7646 21552
rect 6502 21532 7646 21546
rect 6448 21527 6477 21530
rect 7643 21526 7646 21532
rect 7672 21526 7675 21552
rect 8287 21526 8290 21552
rect 8316 21550 8319 21552
rect 8316 21547 8340 21550
rect 8316 21530 8317 21547
rect 8334 21530 8340 21547
rect 8316 21527 8340 21530
rect 10703 21547 10732 21550
rect 10703 21530 10709 21547
rect 10726 21546 10732 21547
rect 10771 21546 10774 21552
rect 10726 21532 10774 21546
rect 10726 21530 10732 21532
rect 10703 21527 10732 21530
rect 8316 21526 8319 21527
rect 10771 21526 10774 21532
rect 10800 21526 10803 21552
rect 12335 21526 12338 21552
rect 12364 21546 12367 21552
rect 12482 21546 12496 21566
rect 12934 21564 12940 21566
rect 12957 21564 12963 21581
rect 12934 21561 12963 21564
rect 15648 21581 15677 21584
rect 15648 21564 15654 21581
rect 15671 21580 15677 21581
rect 19465 21580 19468 21586
rect 15671 21566 19468 21580
rect 15671 21564 15677 21566
rect 15648 21561 15677 21564
rect 19465 21560 19468 21566
rect 19494 21560 19497 21586
rect 29722 21580 29736 21624
rect 29769 21580 29772 21586
rect 29722 21566 29772 21580
rect 29769 21560 29772 21566
rect 29798 21560 29801 21586
rect 12364 21532 12496 21546
rect 12364 21526 12367 21532
rect 12611 21526 12614 21552
rect 12640 21546 12643 21552
rect 12681 21547 12710 21550
rect 12681 21546 12687 21547
rect 12640 21532 12687 21546
rect 12640 21526 12643 21532
rect 12681 21530 12687 21532
rect 12704 21530 12710 21547
rect 12681 21527 12710 21530
rect 29309 21526 29312 21552
rect 29338 21546 29341 21552
rect 29494 21547 29523 21550
rect 29494 21546 29500 21547
rect 29338 21532 29500 21546
rect 29338 21526 29341 21532
rect 29494 21530 29500 21532
rect 29517 21530 29523 21547
rect 29494 21527 29523 21530
rect 3036 21464 29992 21512
rect 3687 21424 3690 21450
rect 3716 21444 3719 21450
rect 6333 21445 6362 21448
rect 3716 21430 6217 21444
rect 3716 21424 3719 21430
rect 4883 21390 4886 21416
rect 4912 21390 4915 21416
rect 6203 21410 6217 21430
rect 6333 21428 6339 21445
rect 6356 21444 6362 21445
rect 6631 21444 6634 21450
rect 6356 21430 6634 21444
rect 6356 21428 6362 21430
rect 6333 21425 6362 21428
rect 6631 21424 6634 21430
rect 6660 21424 6663 21450
rect 7643 21424 7646 21450
rect 7672 21444 7675 21450
rect 8104 21445 8133 21448
rect 8104 21444 8110 21445
rect 7672 21430 8110 21444
rect 7672 21424 7675 21430
rect 8104 21428 8110 21430
rect 8127 21428 8133 21445
rect 8517 21444 8520 21450
rect 8104 21425 8133 21428
rect 8250 21430 8520 21444
rect 8250 21410 8264 21430
rect 8517 21424 8520 21430
rect 8546 21424 8549 21450
rect 9299 21444 9302 21450
rect 8572 21430 9302 21444
rect 6203 21396 8264 21410
rect 8287 21390 8290 21416
rect 8316 21390 8319 21416
rect 4792 21377 4821 21380
rect 4792 21360 4798 21377
rect 4815 21376 4821 21377
rect 4892 21376 4906 21390
rect 4815 21362 4906 21376
rect 4815 21360 4821 21362
rect 4792 21357 4821 21360
rect 4929 21356 4932 21382
rect 4958 21376 4961 21382
rect 8296 21376 8310 21390
rect 8572 21376 8586 21430
rect 9299 21424 9302 21430
rect 9328 21424 9331 21450
rect 9691 21445 9720 21448
rect 9691 21428 9697 21445
rect 9714 21444 9720 21445
rect 10173 21444 10176 21450
rect 9714 21430 10176 21444
rect 9714 21428 9720 21430
rect 9691 21425 9720 21428
rect 10173 21424 10176 21430
rect 10202 21424 10205 21450
rect 12979 21444 12982 21450
rect 10826 21430 12982 21444
rect 4958 21362 5320 21376
rect 4958 21356 4961 21362
rect 4856 21343 4885 21346
rect 4856 21326 4862 21343
rect 4879 21342 4885 21343
rect 5067 21342 5070 21348
rect 4879 21328 5070 21342
rect 4879 21326 4885 21328
rect 4856 21323 4885 21326
rect 5067 21322 5070 21328
rect 5096 21322 5099 21348
rect 5306 21346 5320 21362
rect 8204 21362 8310 21376
rect 8325 21362 8586 21376
rect 8618 21362 8724 21376
rect 5298 21343 5327 21346
rect 5298 21326 5304 21343
rect 5321 21342 5327 21343
rect 5343 21342 5346 21348
rect 5321 21328 5346 21342
rect 5321 21326 5327 21328
rect 5298 21323 5327 21326
rect 5343 21322 5346 21328
rect 5372 21322 5375 21348
rect 5459 21343 5488 21346
rect 5459 21326 5465 21343
rect 5482 21342 5488 21343
rect 5573 21342 5576 21348
rect 5482 21328 5576 21342
rect 5482 21326 5488 21328
rect 5459 21323 5488 21326
rect 5573 21322 5576 21328
rect 5602 21342 5605 21348
rect 5711 21342 5714 21348
rect 5602 21328 5714 21342
rect 5602 21322 5605 21328
rect 5711 21322 5714 21328
rect 5740 21322 5743 21348
rect 8204 21346 8218 21362
rect 8104 21343 8133 21346
rect 8104 21326 8110 21343
rect 8127 21326 8133 21343
rect 8104 21323 8133 21326
rect 8181 21343 8218 21346
rect 8181 21326 8187 21343
rect 8204 21328 8218 21343
rect 8204 21326 8210 21328
rect 8181 21323 8210 21326
rect 4653 21288 4656 21314
rect 4682 21288 4685 21314
rect 4745 21288 4748 21314
rect 4774 21288 4777 21314
rect 4791 21288 4794 21314
rect 4820 21288 4823 21314
rect 5527 21312 5530 21314
rect 5509 21309 5530 21312
rect 5509 21292 5515 21309
rect 5509 21289 5530 21292
rect 5527 21288 5530 21289
rect 5556 21288 5559 21314
rect 8112 21308 8126 21323
rect 8241 21322 8244 21348
rect 8270 21346 8273 21348
rect 8325 21347 8339 21362
rect 8319 21346 8339 21347
rect 8270 21343 8294 21346
rect 8270 21326 8271 21343
rect 8288 21326 8294 21343
rect 8270 21323 8294 21326
rect 8311 21343 8340 21346
rect 8311 21326 8317 21343
rect 8334 21326 8340 21343
rect 8416 21343 8445 21346
rect 8311 21323 8340 21326
rect 8365 21333 8394 21336
rect 8270 21322 8273 21323
rect 8365 21316 8371 21333
rect 8388 21331 8394 21333
rect 8388 21316 8402 21331
rect 8416 21326 8422 21343
rect 8439 21342 8445 21343
rect 8618 21342 8632 21362
rect 8439 21328 8632 21342
rect 8439 21326 8445 21328
rect 8416 21323 8445 21326
rect 8655 21322 8658 21348
rect 8684 21322 8687 21348
rect 8710 21342 8724 21362
rect 10826 21348 10840 21430
rect 12979 21424 12982 21430
rect 13008 21424 13011 21450
rect 16613 21424 16616 21450
rect 16642 21424 16645 21450
rect 26181 21424 26184 21450
rect 26210 21444 26213 21450
rect 29815 21444 29818 21450
rect 26210 21430 29818 21444
rect 26210 21424 26213 21430
rect 29815 21424 29818 21430
rect 29844 21424 29847 21450
rect 20385 21414 20388 21416
rect 20363 21411 20388 21414
rect 20363 21394 20369 21411
rect 20386 21394 20388 21411
rect 20363 21391 20388 21394
rect 20385 21390 20388 21391
rect 20414 21390 20417 21416
rect 24387 21390 24390 21416
rect 24416 21410 24419 21416
rect 25537 21410 25540 21416
rect 24416 21396 25540 21410
rect 24416 21390 24419 21396
rect 25537 21390 25540 21396
rect 25566 21390 25569 21416
rect 10864 21377 10893 21380
rect 10864 21360 10870 21377
rect 10887 21376 10893 21377
rect 15211 21377 15240 21380
rect 10887 21362 11484 21376
rect 10887 21360 10893 21362
rect 10864 21357 10893 21360
rect 9069 21342 9072 21348
rect 8710 21328 9072 21342
rect 9069 21322 9072 21328
rect 9098 21322 9101 21348
rect 10587 21322 10590 21348
rect 10616 21322 10619 21348
rect 10633 21322 10636 21348
rect 10662 21322 10665 21348
rect 10771 21322 10774 21348
rect 10800 21322 10803 21348
rect 10817 21322 10820 21348
rect 10846 21322 10849 21348
rect 11047 21322 11050 21348
rect 11076 21342 11079 21348
rect 11415 21342 11418 21348
rect 11076 21328 11418 21342
rect 11076 21322 11079 21328
rect 11415 21322 11418 21328
rect 11444 21322 11447 21348
rect 11470 21342 11484 21362
rect 15211 21360 15217 21377
rect 15234 21376 15240 21377
rect 16245 21376 16248 21382
rect 15234 21362 16248 21376
rect 15234 21360 15240 21362
rect 15211 21357 15240 21360
rect 16245 21356 16248 21362
rect 16274 21356 16277 21382
rect 19327 21356 19330 21382
rect 19356 21356 19359 21382
rect 21213 21376 21216 21382
rect 20210 21362 21216 21376
rect 13071 21342 13074 21348
rect 11470 21328 13074 21342
rect 13071 21322 13074 21328
rect 13100 21322 13103 21348
rect 14175 21322 14178 21348
rect 14204 21322 14207 21348
rect 16384 21343 16413 21346
rect 16384 21326 16390 21343
rect 16407 21342 16413 21343
rect 16705 21342 16708 21348
rect 16407 21328 16708 21342
rect 16407 21326 16413 21328
rect 16384 21323 16413 21326
rect 16705 21322 16708 21328
rect 16734 21322 16737 21348
rect 16844 21343 16873 21346
rect 16844 21326 16850 21343
rect 16867 21342 16873 21343
rect 17395 21342 17398 21348
rect 16867 21328 17398 21342
rect 16867 21326 16873 21328
rect 16844 21323 16873 21326
rect 17395 21322 17398 21328
rect 17424 21322 17427 21348
rect 19489 21343 19518 21346
rect 19489 21342 19495 21343
rect 19382 21328 19495 21342
rect 8365 21313 8402 21316
rect 8112 21294 8172 21308
rect 7275 21254 7278 21280
rect 7304 21274 7307 21280
rect 7459 21274 7462 21280
rect 7304 21260 7462 21274
rect 7304 21254 7307 21260
rect 7459 21254 7462 21260
rect 7488 21274 7491 21280
rect 7965 21274 7968 21280
rect 7488 21260 7968 21274
rect 7488 21254 7491 21260
rect 7965 21254 7968 21260
rect 7994 21254 7997 21280
rect 8158 21274 8172 21294
rect 8333 21274 8336 21280
rect 8158 21260 8336 21274
rect 8333 21254 8336 21260
rect 8362 21254 8365 21280
rect 8388 21274 8402 21313
rect 8885 21312 8888 21314
rect 8816 21309 8845 21312
rect 8816 21308 8822 21309
rect 8710 21294 8822 21308
rect 8710 21280 8724 21294
rect 8816 21292 8822 21294
rect 8839 21292 8845 21309
rect 8816 21289 8845 21292
rect 8867 21309 8888 21312
rect 8867 21292 8873 21309
rect 8867 21289 8888 21292
rect 8885 21288 8888 21289
rect 8914 21288 8917 21314
rect 10726 21309 10755 21312
rect 10726 21292 10732 21309
rect 10749 21308 10755 21309
rect 10863 21308 10866 21314
rect 10749 21294 10866 21308
rect 10749 21292 10755 21294
rect 10726 21289 10755 21292
rect 10863 21288 10866 21294
rect 10892 21288 10895 21314
rect 10955 21288 10958 21314
rect 10984 21308 10987 21314
rect 11461 21308 11464 21314
rect 10984 21294 11464 21308
rect 10984 21288 10987 21294
rect 11461 21288 11464 21294
rect 11490 21308 11493 21314
rect 11645 21312 11648 21314
rect 11576 21309 11605 21312
rect 11576 21308 11582 21309
rect 11490 21294 11582 21308
rect 11490 21288 11493 21294
rect 11576 21292 11582 21294
rect 11599 21292 11605 21309
rect 11576 21289 11605 21292
rect 11627 21309 11648 21312
rect 11627 21292 11633 21309
rect 11627 21289 11648 21292
rect 11645 21288 11648 21289
rect 11674 21288 11677 21314
rect 13761 21288 13764 21314
rect 13790 21308 13793 21314
rect 14221 21308 14224 21314
rect 13790 21294 14224 21308
rect 13790 21288 13793 21294
rect 14221 21288 14224 21294
rect 14250 21308 14253 21314
rect 14405 21312 14408 21314
rect 14336 21309 14365 21312
rect 14336 21308 14342 21309
rect 14250 21294 14342 21308
rect 14250 21288 14253 21294
rect 14336 21292 14342 21294
rect 14359 21292 14365 21309
rect 14336 21289 14365 21292
rect 14387 21309 14408 21312
rect 14387 21292 14393 21309
rect 14387 21289 14408 21292
rect 14405 21288 14408 21289
rect 14434 21288 14437 21314
rect 19281 21288 19284 21314
rect 19310 21308 19313 21314
rect 19382 21308 19396 21328
rect 19489 21326 19495 21328
rect 19512 21342 19518 21343
rect 20210 21342 20224 21362
rect 21213 21356 21216 21362
rect 21242 21376 21245 21382
rect 21627 21376 21630 21382
rect 21242 21362 21630 21376
rect 21242 21356 21245 21362
rect 21627 21356 21630 21362
rect 21656 21356 21659 21382
rect 23697 21356 23700 21382
rect 23726 21376 23729 21382
rect 24479 21376 24482 21382
rect 23726 21362 24482 21376
rect 23726 21356 23729 21362
rect 24479 21356 24482 21362
rect 24508 21356 24511 21382
rect 19512 21328 20224 21342
rect 19512 21326 19518 21328
rect 19489 21323 19518 21326
rect 20339 21322 20342 21348
rect 20368 21342 20371 21348
rect 24617 21342 24620 21348
rect 20368 21328 24620 21342
rect 20368 21322 20371 21328
rect 24617 21322 24620 21328
rect 24646 21322 24649 21348
rect 19557 21312 19560 21314
rect 19310 21294 19396 21308
rect 19539 21309 19560 21312
rect 19310 21288 19313 21294
rect 19539 21292 19545 21309
rect 19539 21289 19560 21292
rect 19557 21288 19560 21289
rect 19586 21288 19589 21314
rect 24755 21308 24758 21314
rect 20348 21294 24758 21308
rect 8609 21274 8612 21280
rect 8388 21260 8612 21274
rect 8609 21254 8612 21260
rect 8638 21254 8641 21280
rect 8701 21254 8704 21280
rect 8730 21254 8733 21280
rect 9667 21254 9670 21280
rect 9696 21274 9699 21280
rect 10311 21274 10314 21280
rect 9696 21260 10314 21274
rect 9696 21254 9699 21260
rect 10311 21254 10314 21260
rect 10340 21274 10343 21280
rect 11047 21274 11050 21280
rect 10340 21260 11050 21274
rect 10340 21254 10343 21260
rect 11047 21254 11050 21260
rect 11076 21254 11079 21280
rect 12451 21275 12480 21278
rect 12451 21258 12457 21275
rect 12474 21274 12480 21275
rect 12519 21274 12522 21280
rect 12474 21260 12522 21274
rect 12474 21258 12480 21260
rect 12451 21255 12480 21258
rect 12519 21254 12522 21260
rect 12548 21254 12551 21280
rect 20109 21254 20112 21280
rect 20138 21274 20141 21280
rect 20348 21274 20362 21294
rect 24755 21288 24758 21294
rect 24784 21288 24787 21314
rect 20138 21260 20362 21274
rect 20138 21254 20141 21260
rect 3036 21192 29992 21240
rect 3549 21152 3552 21178
rect 3578 21152 3581 21178
rect 6493 21152 6496 21178
rect 6522 21152 6525 21178
rect 6548 21158 7206 21172
rect 3181 21118 3184 21144
rect 3210 21138 3213 21144
rect 3558 21138 3572 21152
rect 3733 21142 3736 21144
rect 3715 21139 3736 21142
rect 3210 21124 3618 21138
rect 3210 21118 3213 21124
rect 3411 21084 3414 21110
rect 3440 21104 3443 21110
rect 3504 21105 3533 21108
rect 3504 21104 3510 21105
rect 3440 21090 3510 21104
rect 3440 21084 3443 21090
rect 3504 21088 3510 21090
rect 3527 21104 3533 21105
rect 3549 21104 3552 21110
rect 3527 21090 3552 21104
rect 3527 21088 3533 21090
rect 3504 21085 3533 21088
rect 3549 21084 3552 21090
rect 3578 21084 3581 21110
rect 3604 21104 3618 21124
rect 3715 21122 3721 21139
rect 3715 21119 3736 21122
rect 3733 21118 3736 21119
rect 3762 21118 3765 21144
rect 4745 21118 4748 21144
rect 4774 21138 4777 21144
rect 6548 21138 6562 21158
rect 4774 21124 6562 21138
rect 4774 21118 4777 21124
rect 6585 21118 6588 21144
rect 6614 21138 6617 21144
rect 6632 21139 6661 21142
rect 6632 21138 6638 21139
rect 6614 21124 6638 21138
rect 6614 21118 6617 21124
rect 6632 21122 6638 21124
rect 6655 21138 6661 21139
rect 6769 21138 6772 21144
rect 6655 21124 6772 21138
rect 6655 21122 6661 21124
rect 6632 21119 6661 21122
rect 6769 21118 6772 21124
rect 6798 21118 6801 21144
rect 3665 21105 3694 21108
rect 3665 21104 3671 21105
rect 3604 21090 3671 21104
rect 3665 21088 3671 21090
rect 3688 21104 3694 21105
rect 3917 21104 3920 21110
rect 3688 21090 3920 21104
rect 3688 21088 3694 21090
rect 3665 21085 3694 21088
rect 3917 21084 3920 21090
rect 3946 21084 3949 21110
rect 4539 21105 4568 21108
rect 4539 21088 4545 21105
rect 4562 21104 4568 21105
rect 4792 21105 4821 21108
rect 4792 21104 4798 21105
rect 4562 21090 4798 21104
rect 4562 21088 4568 21090
rect 4539 21085 4568 21088
rect 4792 21088 4798 21090
rect 4815 21088 4821 21105
rect 4792 21085 4821 21088
rect 4884 21105 4913 21108
rect 4884 21088 4890 21105
rect 4907 21088 4913 21105
rect 4884 21085 4913 21088
rect 4892 21070 4906 21085
rect 4929 21084 4932 21110
rect 4958 21084 4961 21110
rect 4994 21105 5023 21108
rect 4994 21088 5000 21105
rect 5017 21104 5023 21105
rect 5205 21104 5208 21110
rect 5017 21090 5208 21104
rect 5017 21088 5023 21090
rect 4994 21085 5023 21088
rect 5205 21084 5208 21090
rect 5234 21104 5237 21110
rect 5803 21104 5806 21110
rect 5234 21090 5806 21104
rect 5234 21084 5237 21090
rect 5803 21084 5806 21090
rect 5832 21084 5835 21110
rect 6494 21105 6523 21108
rect 6494 21088 6500 21105
rect 6517 21088 6523 21105
rect 6494 21085 6523 21088
rect 5113 21070 5116 21076
rect 4892 21056 5116 21070
rect 5113 21050 5116 21056
rect 5142 21050 5145 21076
rect 4792 21037 4821 21040
rect 4792 21020 4798 21037
rect 4815 21036 4821 21037
rect 4837 21036 4840 21042
rect 4815 21022 4840 21036
rect 4815 21020 4821 21022
rect 4792 21017 4821 21020
rect 4837 21016 4840 21022
rect 4866 21016 4869 21042
rect 6502 21002 6516 21085
rect 6539 21084 6542 21110
rect 6568 21084 6571 21110
rect 6677 21084 6680 21110
rect 6706 21084 6709 21110
rect 6724 21105 6753 21108
rect 6724 21088 6730 21105
rect 6747 21104 6753 21105
rect 6815 21104 6818 21110
rect 6747 21090 6818 21104
rect 6747 21088 6753 21090
rect 6724 21085 6753 21088
rect 6815 21084 6818 21090
rect 6844 21084 6847 21110
rect 7192 21104 7206 21158
rect 8287 21152 8290 21178
rect 8316 21176 8319 21178
rect 8316 21173 8340 21176
rect 8316 21156 8317 21173
rect 8334 21156 8340 21173
rect 8316 21153 8340 21156
rect 10565 21173 10594 21176
rect 10565 21156 10571 21173
rect 10588 21172 10594 21173
rect 10633 21172 10636 21178
rect 10588 21158 10636 21172
rect 10588 21156 10594 21158
rect 10565 21153 10594 21156
rect 8316 21152 8319 21153
rect 10633 21152 10636 21158
rect 10662 21152 10665 21178
rect 12335 21152 12338 21178
rect 12364 21172 12367 21178
rect 12382 21173 12411 21176
rect 12382 21172 12388 21173
rect 12364 21158 12388 21172
rect 12364 21152 12367 21158
rect 12382 21156 12388 21158
rect 12405 21156 12411 21173
rect 12657 21172 12660 21178
rect 12382 21153 12411 21156
rect 12603 21158 12660 21172
rect 7229 21118 7232 21144
rect 7258 21138 7261 21144
rect 7505 21142 7508 21144
rect 7436 21139 7465 21142
rect 7436 21138 7442 21139
rect 7258 21124 7442 21138
rect 7258 21118 7261 21124
rect 7436 21122 7442 21124
rect 7459 21122 7465 21139
rect 7436 21119 7465 21122
rect 7487 21139 7508 21142
rect 7487 21122 7493 21139
rect 7487 21119 7508 21122
rect 7505 21118 7508 21119
rect 7534 21118 7537 21144
rect 9759 21142 9762 21144
rect 9741 21139 9762 21142
rect 9741 21122 9747 21139
rect 9741 21119 9762 21122
rect 9759 21118 9762 21119
rect 9788 21118 9791 21144
rect 12603 21119 12617 21158
rect 12657 21152 12660 21158
rect 12686 21152 12689 21178
rect 13071 21152 13074 21178
rect 13100 21172 13103 21178
rect 16245 21172 16248 21178
rect 13100 21158 16248 21172
rect 13100 21152 13103 21158
rect 16245 21152 16248 21158
rect 16274 21172 16277 21178
rect 16383 21172 16386 21178
rect 16274 21158 16386 21172
rect 16274 21152 16277 21158
rect 16383 21152 16386 21158
rect 16412 21152 16415 21178
rect 20385 21152 20388 21178
rect 20414 21152 20417 21178
rect 23881 21152 23884 21178
rect 23910 21172 23913 21178
rect 23910 21158 25537 21172
rect 23910 21152 23913 21158
rect 12666 21124 12818 21138
rect 12666 21119 12680 21124
rect 12595 21116 12624 21119
rect 7919 21104 7922 21110
rect 7192 21090 7922 21104
rect 7919 21084 7922 21090
rect 7948 21084 7951 21110
rect 7965 21084 7968 21110
rect 7994 21104 7997 21110
rect 7994 21090 8678 21104
rect 7994 21084 7997 21090
rect 8664 21076 8678 21090
rect 8701 21084 8704 21110
rect 8730 21104 8733 21110
rect 9691 21105 9720 21108
rect 9691 21104 9697 21105
rect 8730 21090 9697 21104
rect 8730 21084 8733 21090
rect 9691 21088 9697 21090
rect 9714 21104 9720 21105
rect 9805 21104 9808 21110
rect 9714 21090 9808 21104
rect 9714 21088 9720 21090
rect 9691 21085 9720 21088
rect 9805 21084 9808 21090
rect 9834 21104 9837 21110
rect 10955 21104 10958 21110
rect 9834 21090 10958 21104
rect 9834 21084 9837 21090
rect 10955 21084 10958 21090
rect 10984 21084 10987 21110
rect 12381 21084 12384 21110
rect 12410 21084 12413 21110
rect 12427 21084 12430 21110
rect 12456 21108 12459 21110
rect 12456 21105 12468 21108
rect 12462 21088 12468 21105
rect 12456 21085 12468 21088
rect 12456 21084 12459 21085
rect 12519 21084 12522 21110
rect 12548 21108 12551 21110
rect 12548 21105 12569 21108
rect 12563 21088 12569 21105
rect 12595 21099 12601 21116
rect 12618 21099 12624 21116
rect 12595 21096 12624 21099
rect 12643 21116 12680 21119
rect 12643 21099 12649 21116
rect 12666 21100 12680 21116
rect 12694 21105 12723 21108
rect 12666 21099 12672 21100
rect 12643 21096 12672 21099
rect 12548 21085 12569 21088
rect 12694 21088 12700 21105
rect 12717 21098 12723 21105
rect 12749 21098 12752 21110
rect 12717 21088 12752 21098
rect 12694 21085 12752 21088
rect 12548 21084 12551 21085
rect 12702 21084 12752 21085
rect 12778 21084 12781 21110
rect 7275 21050 7278 21076
rect 7304 21050 7307 21076
rect 8655 21050 8658 21076
rect 8684 21070 8687 21076
rect 9530 21071 9559 21074
rect 9530 21070 9536 21071
rect 8684 21056 9536 21070
rect 8684 21050 8687 21056
rect 9530 21054 9536 21056
rect 9553 21054 9559 21071
rect 11553 21070 11556 21076
rect 9530 21051 9559 21054
rect 11033 21056 11556 21070
rect 7919 21002 7922 21008
rect 6502 20988 7922 21002
rect 7919 20982 7922 20988
rect 7948 20982 7951 21008
rect 9538 21002 9552 21051
rect 9667 21002 9670 21008
rect 9538 20988 9670 21002
rect 9667 20982 9670 20988
rect 9696 20982 9699 21008
rect 10219 20982 10222 21008
rect 10248 21002 10251 21008
rect 11033 21002 11047 21056
rect 11553 21050 11556 21056
rect 11582 21050 11585 21076
rect 12611 21050 12614 21076
rect 12640 21070 12643 21076
rect 12804 21070 12818 21124
rect 12979 21118 12982 21144
rect 13008 21138 13011 21144
rect 17257 21138 17260 21144
rect 13008 21124 17260 21138
rect 13008 21118 13011 21124
rect 17257 21118 17260 21124
rect 17286 21138 17289 21144
rect 18223 21138 18226 21144
rect 17286 21124 18226 21138
rect 17286 21118 17289 21124
rect 18223 21118 18226 21124
rect 18252 21118 18255 21144
rect 18545 21142 18548 21144
rect 18527 21139 18548 21142
rect 18527 21122 18533 21139
rect 18527 21119 18548 21122
rect 18545 21118 18548 21119
rect 18574 21118 18577 21144
rect 19351 21139 19380 21142
rect 19351 21122 19357 21139
rect 19374 21138 19380 21139
rect 20339 21138 20342 21144
rect 19374 21124 20178 21138
rect 19374 21122 19380 21124
rect 19351 21119 19380 21122
rect 12933 21084 12936 21110
rect 12962 21104 12965 21110
rect 16567 21104 16570 21110
rect 12962 21090 16570 21104
rect 12962 21084 12965 21090
rect 16567 21084 16570 21090
rect 16596 21104 16599 21110
rect 17211 21104 17214 21110
rect 16596 21090 17214 21104
rect 16596 21084 16599 21090
rect 17211 21084 17214 21090
rect 17240 21084 17243 21110
rect 18477 21105 18506 21108
rect 18477 21088 18483 21105
rect 18500 21104 18506 21105
rect 18500 21090 19304 21104
rect 18500 21088 18506 21090
rect 18477 21085 18506 21088
rect 19290 21076 19304 21090
rect 20109 21084 20112 21110
rect 20138 21084 20141 21110
rect 20164 21108 20178 21124
rect 20331 21119 20342 21138
rect 20317 21118 20342 21119
rect 20368 21118 20371 21144
rect 20317 21116 20346 21118
rect 20164 21105 20196 21108
rect 20164 21090 20173 21105
rect 20167 21088 20173 21090
rect 20190 21088 20196 21105
rect 20167 21085 20196 21088
rect 20247 21084 20250 21110
rect 20276 21108 20279 21110
rect 20276 21105 20290 21108
rect 20284 21088 20290 21105
rect 20317 21099 20323 21116
rect 20340 21099 20346 21116
rect 20394 21104 20408 21152
rect 20477 21118 20480 21144
rect 20506 21138 20509 21144
rect 23629 21139 23658 21142
rect 23629 21138 23635 21139
rect 20506 21124 23635 21138
rect 20506 21118 20509 21124
rect 23629 21122 23635 21124
rect 23652 21138 23658 21139
rect 25523 21138 25537 21158
rect 26021 21139 26050 21142
rect 26021 21138 26027 21139
rect 23652 21124 23766 21138
rect 25523 21124 26027 21138
rect 23652 21122 23658 21124
rect 23629 21119 23658 21122
rect 20379 21103 20408 21104
rect 20317 21096 20346 21099
rect 20371 21100 20408 21103
rect 20276 21085 20290 21088
rect 20276 21084 20279 21085
rect 20371 21083 20377 21100
rect 20394 21090 20408 21100
rect 20422 21105 20451 21108
rect 20394 21083 20400 21090
rect 20422 21088 20428 21105
rect 20445 21104 20451 21105
rect 20937 21104 20940 21110
rect 20445 21090 20940 21104
rect 20445 21088 20451 21090
rect 20422 21085 20451 21088
rect 20937 21084 20940 21090
rect 20966 21084 20969 21110
rect 23583 21105 23612 21108
rect 23583 21088 23589 21105
rect 23606 21104 23612 21105
rect 23697 21104 23700 21110
rect 23606 21090 23700 21104
rect 23606 21088 23612 21090
rect 23583 21085 23612 21088
rect 23697 21084 23700 21090
rect 23726 21084 23729 21110
rect 23752 21104 23766 21124
rect 26021 21122 26027 21124
rect 26044 21122 26050 21139
rect 26021 21119 26050 21122
rect 23752 21090 25238 21104
rect 20371 21080 20400 21083
rect 12640 21056 12818 21070
rect 12640 21050 12643 21056
rect 14267 21050 14270 21076
rect 14296 21070 14299 21076
rect 14405 21070 14408 21076
rect 14296 21056 14408 21070
rect 14296 21050 14299 21056
rect 14405 21050 14408 21056
rect 14434 21050 14437 21076
rect 18316 21071 18345 21074
rect 18316 21054 18322 21071
rect 18339 21054 18345 21071
rect 18316 21051 18345 21054
rect 12657 21016 12660 21042
rect 12686 21036 12689 21042
rect 16337 21036 16340 21042
rect 12686 21022 16340 21036
rect 12686 21016 12689 21022
rect 16337 21016 16340 21022
rect 16366 21036 16369 21042
rect 17165 21036 17168 21042
rect 16366 21022 17168 21036
rect 16366 21016 16369 21022
rect 17165 21016 17168 21022
rect 17194 21016 17197 21042
rect 10248 20988 11047 21002
rect 18324 21002 18338 21051
rect 19281 21050 19284 21076
rect 19310 21050 19313 21076
rect 23375 21050 23378 21076
rect 23404 21070 23407 21076
rect 23422 21071 23451 21074
rect 23422 21070 23428 21071
rect 23404 21056 23428 21070
rect 23404 21050 23407 21056
rect 23422 21054 23428 21056
rect 23445 21054 23451 21071
rect 23422 21051 23451 21054
rect 19235 21016 19238 21042
rect 19264 21036 19267 21042
rect 20385 21036 20388 21042
rect 19264 21022 20388 21036
rect 19264 21016 19267 21022
rect 20385 21016 20388 21022
rect 20414 21016 20417 21042
rect 20431 21016 20434 21042
rect 20460 21036 20463 21042
rect 20460 21022 23444 21036
rect 20460 21016 20463 21022
rect 19005 21002 19008 21008
rect 18324 20988 19008 21002
rect 10248 20982 10251 20988
rect 19005 20982 19008 20988
rect 19034 21002 19037 21008
rect 19327 21002 19330 21008
rect 19034 20988 19330 21002
rect 19034 20982 19037 20988
rect 19327 20982 19330 20988
rect 19356 20982 19359 21008
rect 20110 21003 20139 21006
rect 20110 20986 20116 21003
rect 20133 21002 20139 21003
rect 22639 21002 22642 21008
rect 20133 20988 22642 21002
rect 20133 20986 20139 20988
rect 20110 20983 20139 20986
rect 22639 20982 22642 20988
rect 22668 20982 22671 21008
rect 23430 21002 23444 21022
rect 23881 21002 23884 21008
rect 23430 20988 23884 21002
rect 23881 20982 23884 20988
rect 23910 20982 23913 21008
rect 24457 21003 24486 21006
rect 24457 20986 24463 21003
rect 24480 21002 24486 21003
rect 24571 21002 24574 21008
rect 24480 20988 24574 21002
rect 24480 20986 24486 20988
rect 24457 20983 24486 20986
rect 24571 20982 24574 20988
rect 24600 20982 24603 21008
rect 25224 21002 25238 21090
rect 25537 21084 25540 21110
rect 25566 21104 25569 21110
rect 25814 21105 25843 21108
rect 25814 21104 25820 21105
rect 25566 21090 25820 21104
rect 25566 21084 25569 21090
rect 25814 21088 25820 21090
rect 25837 21088 25843 21105
rect 25975 21105 26004 21108
rect 25975 21104 25981 21105
rect 25814 21085 25843 21088
rect 25868 21090 25981 21104
rect 25721 21050 25724 21076
rect 25750 21070 25753 21076
rect 25868 21070 25882 21090
rect 25975 21088 25981 21090
rect 25998 21104 26004 21105
rect 26871 21104 26874 21110
rect 25998 21090 26874 21104
rect 25998 21088 26004 21090
rect 25975 21085 26004 21088
rect 26871 21084 26874 21090
rect 26900 21084 26903 21110
rect 25750 21056 25882 21070
rect 25750 21050 25753 21056
rect 26365 21002 26368 21008
rect 25224 20988 26368 21002
rect 26365 20982 26368 20988
rect 26394 20982 26397 21008
rect 26849 21003 26878 21006
rect 26849 20986 26855 21003
rect 26872 21002 26878 21003
rect 27009 21002 27012 21008
rect 26872 20988 27012 21002
rect 26872 20986 26878 20988
rect 26849 20983 26878 20986
rect 27009 20982 27012 20988
rect 27038 20982 27041 21008
rect 3036 20920 29992 20968
rect 3411 20880 3414 20906
rect 3440 20900 3443 20906
rect 4171 20901 4200 20904
rect 3440 20886 4032 20900
rect 3440 20880 3443 20886
rect 4018 20832 4032 20886
rect 4171 20884 4177 20901
rect 4194 20900 4200 20901
rect 4653 20900 4656 20906
rect 4194 20886 4656 20900
rect 4194 20884 4200 20886
rect 4171 20881 4200 20884
rect 4653 20880 4656 20886
rect 4682 20880 4685 20906
rect 6563 20901 6592 20904
rect 6563 20884 6569 20901
rect 6586 20900 6592 20901
rect 6677 20900 6680 20906
rect 6586 20886 6680 20900
rect 6586 20884 6592 20886
rect 6563 20881 6592 20884
rect 6677 20880 6680 20886
rect 6706 20880 6709 20906
rect 7505 20880 7508 20906
rect 7534 20900 7537 20906
rect 7534 20886 8586 20900
rect 7534 20880 7537 20886
rect 6953 20832 6956 20838
rect 4018 20818 5596 20832
rect 3136 20799 3165 20802
rect 3136 20782 3142 20799
rect 3159 20798 3165 20799
rect 3549 20798 3552 20804
rect 3159 20784 3552 20798
rect 3159 20782 3165 20784
rect 3136 20779 3165 20782
rect 3549 20778 3552 20784
rect 3578 20778 3581 20804
rect 5343 20778 5346 20804
rect 5372 20798 5375 20804
rect 5528 20799 5557 20802
rect 5528 20798 5534 20799
rect 5372 20784 5534 20798
rect 5372 20778 5375 20784
rect 5528 20782 5534 20784
rect 5551 20782 5557 20799
rect 5582 20798 5596 20818
rect 6686 20818 6956 20832
rect 6686 20798 6700 20818
rect 6953 20812 6956 20818
rect 6982 20812 6985 20838
rect 7459 20812 7462 20838
rect 7488 20832 7491 20838
rect 7598 20833 7627 20836
rect 7598 20832 7604 20833
rect 7488 20818 7604 20832
rect 7488 20812 7491 20818
rect 7598 20816 7604 20818
rect 7621 20816 7627 20833
rect 7598 20813 7627 20816
rect 5582 20784 6700 20798
rect 5528 20779 5557 20782
rect 6723 20778 6726 20804
rect 6752 20798 6755 20804
rect 6815 20798 6818 20804
rect 6752 20784 6818 20798
rect 6752 20778 6755 20784
rect 6815 20778 6818 20784
rect 6844 20778 6847 20804
rect 7551 20778 7554 20804
rect 7580 20798 7583 20804
rect 7797 20799 7826 20802
rect 7797 20798 7803 20799
rect 7580 20784 7803 20798
rect 7580 20778 7583 20784
rect 7797 20782 7803 20784
rect 7820 20782 7826 20799
rect 8572 20798 8586 20886
rect 8609 20880 8612 20906
rect 8638 20904 8641 20906
rect 8638 20901 8662 20904
rect 8638 20884 8639 20901
rect 8656 20884 8662 20901
rect 8638 20881 8662 20884
rect 8638 20880 8641 20881
rect 9575 20880 9578 20906
rect 9604 20900 9607 20906
rect 11231 20900 11234 20906
rect 9604 20886 11234 20900
rect 9604 20880 9607 20886
rect 11231 20880 11234 20886
rect 11260 20880 11263 20906
rect 11277 20880 11280 20906
rect 11306 20900 11309 20906
rect 11645 20900 11648 20906
rect 11306 20886 11648 20900
rect 11306 20880 11309 20886
rect 11645 20880 11648 20886
rect 11674 20900 11677 20906
rect 13071 20900 13074 20906
rect 11674 20886 13074 20900
rect 11674 20880 11677 20886
rect 13071 20880 13074 20886
rect 13100 20880 13103 20906
rect 14175 20900 14178 20906
rect 13494 20886 14178 20900
rect 12565 20846 12568 20872
rect 12594 20866 12597 20872
rect 12795 20866 12798 20872
rect 12594 20852 12798 20866
rect 12594 20846 12597 20852
rect 12795 20846 12798 20852
rect 12824 20846 12827 20872
rect 10311 20812 10314 20838
rect 10340 20832 10343 20838
rect 10818 20833 10847 20836
rect 10818 20832 10824 20833
rect 10340 20818 10824 20832
rect 10340 20812 10343 20818
rect 10818 20816 10824 20818
rect 10841 20816 10847 20833
rect 10818 20813 10847 20816
rect 11792 20818 11944 20832
rect 8572 20784 8770 20798
rect 7797 20779 7826 20782
rect 3181 20744 3184 20770
rect 3210 20764 3213 20770
rect 3296 20765 3325 20768
rect 3296 20764 3302 20765
rect 3210 20750 3302 20764
rect 3210 20744 3213 20750
rect 3296 20748 3302 20750
rect 3319 20748 3325 20765
rect 3296 20745 3325 20748
rect 3347 20765 3376 20768
rect 3347 20748 3353 20765
rect 3370 20764 3376 20765
rect 3411 20764 3414 20770
rect 3370 20750 3414 20764
rect 3370 20748 3376 20750
rect 3347 20745 3376 20748
rect 3411 20744 3414 20750
rect 3440 20744 3443 20770
rect 5757 20768 5760 20770
rect 5688 20765 5717 20768
rect 5688 20764 5694 20765
rect 5536 20750 5694 20764
rect 5536 20736 5550 20750
rect 5688 20748 5694 20750
rect 5711 20748 5717 20765
rect 5688 20745 5717 20748
rect 5739 20765 5760 20768
rect 5739 20748 5745 20765
rect 5739 20745 5760 20748
rect 5757 20744 5760 20745
rect 5786 20744 5789 20770
rect 7758 20765 7787 20768
rect 7758 20764 7764 20765
rect 7652 20750 7764 20764
rect 3917 20710 3920 20736
rect 3946 20730 3949 20736
rect 5527 20730 5530 20736
rect 3946 20716 5530 20730
rect 3946 20710 3949 20716
rect 5527 20710 5530 20716
rect 5556 20710 5559 20736
rect 6355 20710 6358 20736
rect 6384 20730 6387 20736
rect 7229 20730 7232 20736
rect 6384 20716 7232 20730
rect 6384 20710 6387 20716
rect 7229 20710 7232 20716
rect 7258 20730 7261 20736
rect 7652 20730 7666 20750
rect 7758 20748 7764 20750
rect 7781 20748 7787 20765
rect 8756 20764 8770 20784
rect 10955 20778 10958 20804
rect 10984 20802 10987 20804
rect 10984 20799 11002 20802
rect 10996 20782 11002 20799
rect 10984 20779 11002 20782
rect 11017 20799 11046 20802
rect 11017 20782 11023 20799
rect 11040 20798 11046 20799
rect 11792 20798 11806 20818
rect 11040 20784 11806 20798
rect 11040 20782 11047 20784
rect 11017 20779 11047 20782
rect 10984 20778 10987 20779
rect 11033 20764 11047 20779
rect 11829 20778 11832 20804
rect 11858 20802 11861 20804
rect 11858 20799 11882 20802
rect 11858 20782 11859 20799
rect 11876 20782 11882 20799
rect 11930 20798 11944 20818
rect 12933 20812 12936 20838
rect 12962 20832 12965 20838
rect 13494 20836 13508 20886
rect 14175 20880 14178 20886
rect 14204 20880 14207 20906
rect 17993 20880 17996 20906
rect 18022 20900 18025 20906
rect 18545 20900 18548 20906
rect 18022 20886 18548 20900
rect 18022 20880 18025 20886
rect 18545 20880 18548 20886
rect 18574 20900 18577 20906
rect 20041 20901 20070 20904
rect 18574 20886 19856 20900
rect 18574 20880 18577 20886
rect 19842 20866 19856 20886
rect 20041 20884 20047 20901
rect 20064 20900 20070 20901
rect 20247 20900 20250 20906
rect 20064 20886 20250 20900
rect 20064 20884 20070 20886
rect 20041 20881 20070 20884
rect 20247 20880 20250 20886
rect 20276 20880 20279 20906
rect 28067 20900 28070 20906
rect 27984 20886 28070 20900
rect 20431 20866 20434 20872
rect 19842 20852 20434 20866
rect 20431 20846 20434 20852
rect 20460 20846 20463 20872
rect 13486 20833 13515 20836
rect 13486 20832 13492 20833
rect 12962 20818 13492 20832
rect 12962 20812 12965 20818
rect 13486 20816 13492 20818
rect 13509 20816 13515 20833
rect 13486 20813 13515 20816
rect 19005 20812 19008 20838
rect 19034 20812 19037 20838
rect 22501 20812 22504 20838
rect 22530 20812 22533 20838
rect 24663 20812 24666 20838
rect 24692 20812 24695 20838
rect 26871 20812 26874 20838
rect 26900 20832 26903 20838
rect 27984 20836 27998 20886
rect 28067 20880 28070 20886
rect 28096 20900 28099 20906
rect 28205 20900 28208 20906
rect 28096 20886 28208 20900
rect 28096 20880 28099 20886
rect 28205 20880 28208 20886
rect 28234 20880 28237 20906
rect 27976 20833 28005 20836
rect 26900 20818 27124 20832
rect 26900 20812 26903 20818
rect 13301 20798 13304 20804
rect 11930 20784 13304 20798
rect 11858 20779 11882 20782
rect 11858 20778 11861 20779
rect 13301 20778 13304 20784
rect 13330 20778 13333 20804
rect 13685 20799 13714 20802
rect 13685 20798 13691 20799
rect 13494 20784 13691 20798
rect 8756 20750 11047 20764
rect 7758 20745 7787 20748
rect 13025 20744 13028 20770
rect 13054 20764 13057 20770
rect 13494 20764 13508 20784
rect 13685 20782 13691 20784
rect 13708 20782 13714 20799
rect 13685 20779 13714 20782
rect 19167 20799 19196 20802
rect 19167 20782 19173 20799
rect 19190 20798 19196 20799
rect 19281 20798 19284 20804
rect 19190 20784 19284 20798
rect 19190 20782 19196 20784
rect 19167 20779 19196 20782
rect 19281 20778 19284 20784
rect 19310 20778 19313 20804
rect 21075 20778 21078 20804
rect 21104 20798 21107 20804
rect 21214 20799 21243 20802
rect 21214 20798 21220 20799
rect 21104 20784 21220 20798
rect 21104 20778 21107 20784
rect 21214 20782 21220 20784
rect 21237 20782 21243 20799
rect 21214 20779 21243 20782
rect 22639 20778 22642 20804
rect 22668 20778 22671 20804
rect 24755 20778 24758 20804
rect 24784 20802 24787 20804
rect 24784 20798 24788 20802
rect 27055 20798 27058 20804
rect 24784 20784 27058 20798
rect 24784 20779 24788 20784
rect 24784 20778 24787 20779
rect 27055 20778 27058 20784
rect 27084 20778 27087 20804
rect 27110 20798 27124 20818
rect 27976 20816 27982 20833
rect 27999 20816 28005 20833
rect 27976 20813 28005 20816
rect 28113 20798 28116 20804
rect 28142 20802 28145 20804
rect 28142 20799 28160 20802
rect 27110 20784 28116 20798
rect 28113 20778 28116 20784
rect 28154 20782 28160 20799
rect 28142 20779 28160 20782
rect 28175 20799 28204 20802
rect 28175 20782 28181 20799
rect 28198 20798 28204 20799
rect 28251 20798 28254 20804
rect 28198 20784 28254 20798
rect 28198 20782 28204 20784
rect 28175 20779 28204 20782
rect 28142 20778 28145 20779
rect 28251 20778 28254 20784
rect 28280 20778 28283 20804
rect 13646 20765 13675 20768
rect 13646 20764 13652 20765
rect 13054 20750 13508 20764
rect 13540 20750 13652 20764
rect 13054 20744 13057 20750
rect 7258 20716 7666 20730
rect 7258 20710 7261 20716
rect 11277 20710 11280 20736
rect 11306 20730 11309 20736
rect 12611 20730 12614 20736
rect 11306 20716 12614 20730
rect 11306 20710 11309 20716
rect 12611 20710 12614 20716
rect 12640 20730 12643 20736
rect 13071 20730 13074 20736
rect 12640 20716 13074 20730
rect 12640 20710 12643 20716
rect 13071 20710 13074 20716
rect 13100 20730 13103 20736
rect 13540 20730 13554 20750
rect 13646 20748 13652 20750
rect 13669 20764 13675 20765
rect 13761 20764 13764 20770
rect 13669 20750 13764 20764
rect 13669 20748 13675 20750
rect 13646 20745 13675 20748
rect 13761 20744 13764 20750
rect 13790 20744 13793 20770
rect 19235 20768 19238 20770
rect 19217 20765 19238 20768
rect 19217 20748 19223 20765
rect 19217 20745 19238 20748
rect 19235 20744 19238 20745
rect 19264 20744 19267 20770
rect 21443 20768 21446 20770
rect 21375 20765 21404 20768
rect 21375 20764 21381 20765
rect 21222 20750 21381 20764
rect 21222 20736 21236 20750
rect 21375 20748 21381 20750
rect 21398 20748 21404 20765
rect 21375 20745 21404 20748
rect 21425 20765 21446 20768
rect 21425 20748 21431 20765
rect 21425 20745 21446 20748
rect 21443 20744 21446 20745
rect 21472 20744 21475 20770
rect 22685 20744 22688 20770
rect 22714 20744 22717 20770
rect 22869 20744 22872 20770
rect 22898 20744 22901 20770
rect 24571 20744 24574 20770
rect 24600 20744 24603 20770
rect 24617 20744 24620 20770
rect 24646 20764 24649 20770
rect 24664 20765 24693 20768
rect 24664 20764 24670 20765
rect 24646 20750 24670 20764
rect 24646 20744 24649 20750
rect 24664 20748 24670 20750
rect 24687 20748 24693 20765
rect 24664 20745 24693 20748
rect 13100 20716 13554 20730
rect 14521 20731 14550 20734
rect 13100 20710 13103 20716
rect 14521 20714 14527 20731
rect 14544 20730 14550 20731
rect 14865 20730 14868 20736
rect 14544 20716 14868 20730
rect 14544 20714 14550 20716
rect 14521 20711 14550 20714
rect 14865 20710 14868 20716
rect 14894 20710 14897 20736
rect 21213 20710 21216 20736
rect 21242 20710 21245 20736
rect 22249 20731 22278 20734
rect 22249 20714 22255 20731
rect 22272 20730 22278 20731
rect 22547 20730 22550 20736
rect 22272 20716 22550 20730
rect 22272 20714 22278 20716
rect 22249 20711 22278 20714
rect 22547 20710 22550 20716
rect 22576 20710 22579 20736
rect 22593 20710 22596 20736
rect 22622 20710 22625 20736
rect 24672 20730 24686 20745
rect 24709 20744 24712 20770
rect 24738 20744 24741 20770
rect 27193 20730 27196 20736
rect 24672 20716 27196 20730
rect 27193 20710 27196 20716
rect 27222 20710 27225 20736
rect 29011 20731 29040 20734
rect 29011 20714 29017 20731
rect 29034 20730 29040 20731
rect 29585 20730 29588 20736
rect 29034 20716 29588 20730
rect 29034 20714 29040 20716
rect 29011 20711 29040 20714
rect 29585 20710 29588 20716
rect 29614 20710 29617 20736
rect 3036 20648 29992 20696
rect 4815 20629 4844 20632
rect 4815 20612 4821 20629
rect 4838 20628 4844 20629
rect 4929 20628 4932 20634
rect 4838 20614 4932 20628
rect 4838 20612 4844 20614
rect 4815 20609 4844 20612
rect 4929 20608 4932 20614
rect 4958 20608 4961 20634
rect 5527 20608 5530 20634
rect 5556 20628 5559 20634
rect 5711 20628 5714 20634
rect 5556 20614 5714 20628
rect 5556 20608 5559 20614
rect 5711 20608 5714 20614
rect 5740 20628 5743 20634
rect 5740 20614 6217 20628
rect 5740 20608 5743 20614
rect 3825 20574 3828 20600
rect 3854 20594 3857 20600
rect 3979 20595 4008 20598
rect 3979 20594 3985 20595
rect 3854 20580 3985 20594
rect 3854 20574 3857 20580
rect 3979 20578 3985 20580
rect 4002 20594 4008 20595
rect 6203 20594 6217 20614
rect 7919 20608 7922 20634
rect 7948 20608 7951 20634
rect 15509 20608 15512 20634
rect 15538 20608 15541 20634
rect 24549 20629 24578 20632
rect 24549 20612 24555 20629
rect 24572 20628 24578 20629
rect 24709 20628 24712 20634
rect 24572 20614 24712 20628
rect 24572 20612 24578 20614
rect 24549 20609 24578 20612
rect 24709 20608 24712 20614
rect 24738 20608 24741 20634
rect 29585 20608 29588 20634
rect 29614 20628 29617 20634
rect 29614 20614 29685 20628
rect 29614 20608 29617 20614
rect 6355 20594 6358 20600
rect 4002 20580 4124 20594
rect 6203 20580 6358 20594
rect 4002 20578 4008 20580
rect 3979 20575 4008 20578
rect 3549 20540 3552 20566
rect 3578 20560 3581 20566
rect 3780 20561 3809 20564
rect 3780 20560 3786 20561
rect 3578 20546 3786 20560
rect 3578 20540 3581 20546
rect 3780 20544 3786 20546
rect 3803 20544 3809 20561
rect 3780 20541 3809 20544
rect 3917 20540 3920 20566
rect 3946 20564 3949 20566
rect 3946 20561 3964 20564
rect 3958 20544 3964 20561
rect 4110 20560 4124 20580
rect 6355 20574 6358 20580
rect 6384 20574 6387 20600
rect 7597 20574 7600 20600
rect 7626 20594 7629 20600
rect 7626 20580 7896 20594
rect 7626 20574 7629 20580
rect 4469 20560 4472 20566
rect 4110 20546 4472 20560
rect 3946 20541 3964 20544
rect 3946 20540 3949 20541
rect 4469 20540 4472 20546
rect 4498 20540 4501 20566
rect 6364 20560 6378 20574
rect 6493 20560 6496 20566
rect 6522 20564 6525 20566
rect 6522 20561 6540 20564
rect 6364 20546 6496 20560
rect 6493 20540 6496 20546
rect 6534 20544 6540 20561
rect 6522 20541 6540 20544
rect 6555 20561 6584 20564
rect 6555 20544 6561 20561
rect 6578 20560 6584 20561
rect 6999 20560 7002 20566
rect 6578 20546 7002 20560
rect 6578 20544 6584 20546
rect 6555 20541 6584 20544
rect 6522 20540 6525 20541
rect 6999 20540 7002 20546
rect 7028 20540 7031 20566
rect 7391 20561 7420 20564
rect 7391 20544 7397 20561
rect 7414 20560 7420 20561
rect 7644 20561 7673 20564
rect 7644 20560 7650 20561
rect 7414 20546 7650 20560
rect 7414 20544 7420 20546
rect 7391 20541 7420 20544
rect 7644 20544 7650 20546
rect 7667 20544 7673 20561
rect 7644 20541 7673 20544
rect 7689 20540 7692 20566
rect 7718 20560 7721 20566
rect 7736 20561 7765 20564
rect 7736 20560 7742 20561
rect 7718 20546 7742 20560
rect 7718 20540 7721 20546
rect 7736 20544 7742 20546
rect 7759 20544 7765 20561
rect 7736 20541 7765 20544
rect 7781 20540 7784 20566
rect 7810 20540 7813 20566
rect 7827 20540 7830 20566
rect 7856 20540 7859 20566
rect 7882 20560 7896 20580
rect 9653 20580 11786 20594
rect 8287 20560 8290 20566
rect 7882 20546 8290 20560
rect 8287 20540 8290 20546
rect 8316 20560 8319 20566
rect 9653 20560 9667 20580
rect 8316 20546 9667 20560
rect 8316 20540 8319 20546
rect 11369 20540 11372 20566
rect 11398 20560 11401 20566
rect 11461 20560 11464 20566
rect 11398 20546 11464 20560
rect 11398 20540 11401 20546
rect 11461 20540 11464 20546
rect 11490 20560 11493 20566
rect 11772 20564 11786 20580
rect 14221 20574 14224 20600
rect 14250 20594 14253 20600
rect 15418 20595 15447 20598
rect 15418 20594 15424 20595
rect 14250 20580 15424 20594
rect 14250 20574 14253 20580
rect 15418 20578 15424 20580
rect 15441 20578 15447 20595
rect 15418 20575 15447 20578
rect 21121 20574 21124 20600
rect 21150 20594 21153 20600
rect 21287 20595 21316 20598
rect 21287 20594 21293 20595
rect 21150 20580 21293 20594
rect 21150 20574 21153 20580
rect 21287 20578 21293 20580
rect 21310 20594 21316 20595
rect 21310 20580 21420 20594
rect 21310 20578 21316 20580
rect 21287 20575 21316 20578
rect 11709 20561 11738 20564
rect 11709 20560 11715 20561
rect 11490 20546 11715 20560
rect 11490 20540 11493 20546
rect 11709 20544 11715 20546
rect 11732 20544 11738 20561
rect 11709 20541 11738 20544
rect 11753 20561 11786 20564
rect 11753 20544 11759 20561
rect 11776 20560 11786 20561
rect 11776 20546 12450 20560
rect 11776 20544 11782 20546
rect 11753 20541 11782 20544
rect 6171 20506 6174 20532
rect 6200 20526 6203 20532
rect 6356 20527 6385 20530
rect 6356 20526 6362 20527
rect 6200 20512 6362 20526
rect 6200 20506 6203 20512
rect 6356 20510 6362 20512
rect 6379 20510 6385 20527
rect 7836 20526 7850 20540
rect 10265 20526 10268 20532
rect 6356 20507 6385 20510
rect 7652 20512 10268 20526
rect 7652 20498 7666 20512
rect 10265 20506 10268 20512
rect 10294 20506 10297 20532
rect 11047 20506 11050 20532
rect 11076 20526 11079 20532
rect 11415 20526 11418 20532
rect 11076 20512 11418 20526
rect 11076 20506 11079 20512
rect 11415 20506 11418 20512
rect 11444 20526 11447 20532
rect 11554 20527 11583 20530
rect 11554 20526 11560 20527
rect 11444 20512 11560 20526
rect 11444 20506 11447 20512
rect 11554 20510 11560 20512
rect 11577 20510 11583 20527
rect 11554 20507 11583 20510
rect 7643 20472 7646 20498
rect 7672 20472 7675 20498
rect 7689 20472 7692 20498
rect 7718 20492 7721 20498
rect 8977 20492 8980 20498
rect 7718 20478 8980 20492
rect 7718 20472 7721 20478
rect 8977 20472 8980 20478
rect 9006 20492 9009 20498
rect 10173 20492 10176 20498
rect 9006 20478 10176 20492
rect 9006 20472 9009 20478
rect 10173 20472 10176 20478
rect 10202 20472 10205 20498
rect 12436 20492 12450 20546
rect 14773 20540 14776 20566
rect 14802 20540 14805 20566
rect 14865 20540 14868 20566
rect 14894 20540 14897 20566
rect 15279 20540 15282 20566
rect 15308 20540 15311 20566
rect 15326 20561 15355 20564
rect 15326 20544 15332 20561
rect 15349 20544 15355 20561
rect 15326 20541 15355 20544
rect 12795 20506 12798 20532
rect 12824 20526 12827 20532
rect 13025 20526 13028 20532
rect 12824 20512 13028 20526
rect 12824 20506 12827 20512
rect 13025 20506 13028 20512
rect 13054 20506 13057 20532
rect 14782 20492 14796 20540
rect 14820 20527 14849 20530
rect 14820 20510 14826 20527
rect 14843 20526 14849 20527
rect 15334 20526 15348 20541
rect 15371 20540 15374 20566
rect 15400 20540 15403 20566
rect 21213 20540 21216 20566
rect 21242 20564 21245 20566
rect 21242 20561 21266 20564
rect 21242 20544 21243 20561
rect 21260 20560 21266 20561
rect 21351 20560 21354 20566
rect 21260 20546 21354 20560
rect 21260 20544 21266 20546
rect 21242 20541 21266 20544
rect 21242 20540 21245 20541
rect 21351 20540 21354 20546
rect 21380 20540 21383 20566
rect 21406 20560 21420 20580
rect 22547 20574 22550 20600
rect 22576 20594 22579 20600
rect 22594 20595 22623 20598
rect 22594 20594 22600 20595
rect 22576 20580 22600 20594
rect 22576 20574 22579 20580
rect 22594 20578 22600 20580
rect 22617 20578 22623 20595
rect 22594 20575 22623 20578
rect 23725 20595 23754 20598
rect 23725 20578 23731 20595
rect 23748 20594 23754 20595
rect 23748 20580 23858 20594
rect 23748 20578 23754 20580
rect 23725 20575 23754 20578
rect 21406 20546 22064 20560
rect 14843 20512 15348 20526
rect 14843 20510 14849 20512
rect 14820 20507 14849 20510
rect 21075 20506 21078 20532
rect 21104 20506 21107 20532
rect 15003 20492 15006 20498
rect 12436 20478 13048 20492
rect 14782 20478 15006 20492
rect 13034 20464 13048 20478
rect 15003 20472 15006 20478
rect 15032 20472 15035 20498
rect 12381 20438 12384 20464
rect 12410 20458 12413 20464
rect 12589 20459 12618 20462
rect 12589 20458 12595 20459
rect 12410 20444 12595 20458
rect 12410 20438 12413 20444
rect 12589 20442 12595 20444
rect 12612 20442 12618 20459
rect 12589 20439 12618 20442
rect 13025 20438 13028 20464
rect 13054 20458 13057 20464
rect 13439 20458 13442 20464
rect 13054 20444 13442 20458
rect 13054 20438 13057 20444
rect 13439 20438 13442 20444
rect 13468 20438 13471 20464
rect 15923 20438 15926 20464
rect 15952 20458 15955 20464
rect 17027 20458 17030 20464
rect 15952 20444 17030 20458
rect 15952 20438 15955 20444
rect 17027 20438 17030 20444
rect 17056 20438 17059 20464
rect 22050 20458 22064 20546
rect 22639 20540 22642 20566
rect 22668 20560 22671 20566
rect 22686 20561 22715 20564
rect 22686 20560 22692 20561
rect 22668 20546 22692 20560
rect 22668 20540 22671 20546
rect 22686 20544 22692 20546
rect 22709 20544 22715 20561
rect 22686 20541 22715 20544
rect 22732 20561 22761 20564
rect 22732 20544 22738 20561
rect 22755 20544 22761 20561
rect 22732 20541 22761 20544
rect 22796 20561 22825 20564
rect 22796 20544 22802 20561
rect 22819 20560 22825 20561
rect 22915 20560 22918 20566
rect 22819 20546 22918 20560
rect 22819 20544 22825 20546
rect 22796 20541 22825 20544
rect 22111 20527 22140 20530
rect 22111 20510 22117 20527
rect 22134 20526 22140 20527
rect 22740 20526 22754 20541
rect 22915 20540 22918 20546
rect 22944 20540 22947 20566
rect 23559 20540 23562 20566
rect 23588 20560 23591 20566
rect 23651 20560 23654 20566
rect 23680 20564 23683 20566
rect 23680 20561 23698 20564
rect 23588 20546 23654 20560
rect 23588 20540 23591 20546
rect 23651 20540 23654 20546
rect 23692 20544 23698 20561
rect 23844 20560 23858 20580
rect 25583 20574 25586 20600
rect 25612 20594 25615 20600
rect 25737 20595 25766 20598
rect 25737 20594 25743 20595
rect 25612 20580 25743 20594
rect 25612 20574 25615 20580
rect 25737 20578 25743 20580
rect 25760 20578 25766 20595
rect 25737 20575 25766 20578
rect 28113 20574 28116 20600
rect 28142 20594 28145 20600
rect 28274 20595 28303 20598
rect 28274 20594 28280 20595
rect 28142 20580 28280 20594
rect 28142 20574 28145 20580
rect 28274 20578 28280 20580
rect 28297 20578 28303 20595
rect 28274 20575 28303 20578
rect 29149 20595 29178 20598
rect 29149 20578 29155 20595
rect 29172 20594 29178 20595
rect 29172 20580 29470 20594
rect 29172 20578 29178 20580
rect 29149 20575 29178 20578
rect 23927 20560 23930 20566
rect 23844 20546 23930 20560
rect 23680 20541 23698 20544
rect 23680 20540 23683 20541
rect 23927 20540 23930 20546
rect 23956 20540 23959 20566
rect 25675 20540 25678 20566
rect 25704 20564 25707 20566
rect 25704 20561 25722 20564
rect 25716 20544 25722 20561
rect 25704 20541 25722 20544
rect 25704 20540 25707 20541
rect 26825 20540 26828 20566
rect 26854 20540 26857 20566
rect 26918 20561 26947 20564
rect 26918 20544 26924 20561
rect 26941 20544 26947 20561
rect 26918 20541 26947 20544
rect 28313 20561 28342 20564
rect 28313 20544 28319 20561
rect 28336 20560 28342 20561
rect 28527 20560 28530 20566
rect 28336 20546 28530 20560
rect 28336 20544 28342 20546
rect 28313 20541 28342 20544
rect 22134 20512 22754 20526
rect 22134 20510 22140 20512
rect 22111 20507 22140 20510
rect 23053 20506 23056 20532
rect 23082 20526 23085 20532
rect 23375 20526 23378 20532
rect 23082 20512 23378 20526
rect 23082 20506 23085 20512
rect 23375 20506 23378 20512
rect 23404 20526 23407 20532
rect 23514 20527 23543 20530
rect 23514 20526 23520 20527
rect 23404 20512 23520 20526
rect 23404 20506 23407 20512
rect 23514 20510 23520 20512
rect 23537 20510 23543 20527
rect 23514 20507 23543 20510
rect 25537 20506 25540 20532
rect 25566 20506 25569 20532
rect 22594 20493 22623 20496
rect 22594 20476 22600 20493
rect 22617 20492 22623 20493
rect 22685 20492 22688 20498
rect 22617 20478 22688 20492
rect 22617 20476 22623 20478
rect 22594 20473 22623 20476
rect 22685 20472 22688 20478
rect 22714 20472 22717 20498
rect 26872 20493 26901 20496
rect 26872 20492 26878 20493
rect 26374 20478 26878 20492
rect 23237 20458 23240 20464
rect 22050 20444 23240 20458
rect 23237 20438 23240 20444
rect 23266 20438 23269 20464
rect 26227 20438 26230 20464
rect 26256 20458 26259 20464
rect 26374 20458 26388 20478
rect 26872 20476 26878 20478
rect 26895 20476 26901 20493
rect 26872 20473 26901 20476
rect 26256 20444 26388 20458
rect 26573 20459 26602 20462
rect 26256 20438 26259 20444
rect 26573 20442 26579 20459
rect 26596 20458 26602 20459
rect 26779 20458 26782 20464
rect 26596 20444 26782 20458
rect 26596 20442 26602 20444
rect 26573 20439 26602 20442
rect 26779 20438 26782 20444
rect 26808 20438 26811 20464
rect 26926 20458 26940 20541
rect 28527 20540 28530 20546
rect 28556 20540 28559 20566
rect 29355 20540 29358 20566
rect 29384 20560 29387 20566
rect 29456 20564 29470 20580
rect 29671 20567 29685 20614
rect 29402 20561 29431 20564
rect 29402 20560 29408 20561
rect 29384 20546 29408 20560
rect 29384 20540 29387 20546
rect 29402 20544 29408 20546
rect 29425 20544 29431 20561
rect 29456 20561 29488 20564
rect 29456 20546 29465 20561
rect 29402 20541 29431 20544
rect 29459 20544 29465 20546
rect 29482 20544 29488 20561
rect 29459 20541 29488 20544
rect 29539 20540 29542 20566
rect 29568 20564 29571 20566
rect 29663 20564 29692 20567
rect 29568 20561 29582 20564
rect 29576 20544 29582 20561
rect 29568 20541 29582 20544
rect 29615 20561 29644 20564
rect 29615 20544 29621 20561
rect 29638 20544 29644 20561
rect 29663 20547 29669 20564
rect 29686 20547 29692 20564
rect 29663 20544 29692 20547
rect 29714 20561 29743 20564
rect 29714 20544 29720 20561
rect 29737 20560 29743 20561
rect 29815 20560 29818 20566
rect 29737 20546 29818 20560
rect 29737 20544 29743 20546
rect 29615 20541 29644 20544
rect 29714 20541 29743 20544
rect 29568 20540 29571 20541
rect 28067 20506 28070 20532
rect 28096 20526 28099 20532
rect 28114 20527 28143 20530
rect 28114 20526 28120 20527
rect 28096 20512 28120 20526
rect 28096 20506 28099 20512
rect 28114 20510 28120 20512
rect 28137 20510 28143 20527
rect 28114 20507 28143 20510
rect 29263 20506 29266 20532
rect 29292 20526 29295 20532
rect 29623 20526 29637 20541
rect 29815 20540 29818 20546
rect 29844 20540 29847 20566
rect 29769 20526 29772 20532
rect 29292 20512 29772 20526
rect 29292 20506 29295 20512
rect 29769 20506 29772 20512
rect 29798 20506 29801 20532
rect 29402 20459 29431 20462
rect 29402 20458 29408 20459
rect 26926 20444 29408 20458
rect 29402 20442 29408 20444
rect 29425 20442 29431 20459
rect 29402 20439 29431 20442
rect 3036 20376 29992 20424
rect 5527 20356 5530 20362
rect 5352 20342 5530 20356
rect 5352 20288 5366 20342
rect 5527 20336 5530 20342
rect 5556 20336 5559 20362
rect 6379 20357 6408 20360
rect 6379 20340 6385 20357
rect 6402 20356 6408 20357
rect 6539 20356 6542 20362
rect 6402 20342 6542 20356
rect 6402 20340 6408 20342
rect 6379 20337 6408 20340
rect 6539 20336 6542 20342
rect 6568 20336 6571 20362
rect 9023 20336 9026 20362
rect 9052 20356 9055 20362
rect 11875 20356 11878 20362
rect 9052 20342 11878 20356
rect 9052 20336 9055 20342
rect 11875 20336 11878 20342
rect 11904 20336 11907 20362
rect 12013 20336 12016 20362
rect 12042 20356 12045 20362
rect 12749 20356 12752 20362
rect 12042 20342 12752 20356
rect 12042 20336 12045 20342
rect 12749 20336 12752 20342
rect 12778 20356 12781 20362
rect 12778 20342 13784 20356
rect 12778 20336 12781 20342
rect 13770 20322 13784 20342
rect 14221 20336 14224 20362
rect 14250 20336 14253 20362
rect 15371 20336 15374 20362
rect 15400 20356 15403 20362
rect 17258 20357 17287 20360
rect 17258 20356 17264 20357
rect 15400 20342 17264 20356
rect 15400 20336 15403 20342
rect 17258 20340 17264 20342
rect 17281 20340 17287 20357
rect 17258 20337 17287 20340
rect 19373 20336 19376 20362
rect 19402 20356 19405 20362
rect 19787 20356 19790 20362
rect 19402 20342 19790 20356
rect 19402 20336 19405 20342
rect 19787 20336 19790 20342
rect 19816 20336 19819 20362
rect 21443 20336 21446 20362
rect 21472 20356 21475 20362
rect 25583 20356 25586 20362
rect 21472 20342 25586 20356
rect 21472 20336 21475 20342
rect 25583 20336 25586 20342
rect 25612 20336 25615 20362
rect 26734 20357 26763 20360
rect 26734 20340 26740 20357
rect 26757 20356 26763 20357
rect 26825 20356 26828 20362
rect 26757 20342 26828 20356
rect 26757 20340 26763 20342
rect 26734 20337 26763 20340
rect 26825 20336 26828 20342
rect 26854 20336 26857 20362
rect 28251 20336 28254 20362
rect 28280 20356 28283 20362
rect 28435 20356 28438 20362
rect 28280 20342 28438 20356
rect 28280 20336 28283 20342
rect 28435 20336 28438 20342
rect 28464 20336 28467 20362
rect 29011 20357 29040 20360
rect 29011 20340 29017 20357
rect 29034 20356 29040 20357
rect 29539 20356 29542 20362
rect 29034 20342 29542 20356
rect 29034 20340 29040 20342
rect 29011 20337 29040 20340
rect 29539 20336 29542 20342
rect 29568 20336 29571 20362
rect 13770 20308 15164 20322
rect 5352 20274 5412 20288
rect 3549 20234 3552 20260
rect 3578 20254 3581 20260
rect 5343 20254 5346 20260
rect 3578 20240 5346 20254
rect 3578 20234 3581 20240
rect 5343 20234 5346 20240
rect 5372 20234 5375 20260
rect 5398 20254 5412 20274
rect 11415 20268 11418 20294
rect 11444 20268 11447 20294
rect 12749 20268 12752 20294
rect 12778 20288 12781 20294
rect 12933 20288 12936 20294
rect 12778 20274 12936 20288
rect 12778 20268 12781 20274
rect 12933 20268 12936 20274
rect 12962 20268 12965 20294
rect 5505 20255 5534 20258
rect 5505 20254 5511 20255
rect 5398 20240 5511 20254
rect 5505 20238 5511 20240
rect 5528 20238 5534 20255
rect 5757 20254 5760 20260
rect 5505 20235 5534 20238
rect 5674 20240 5760 20254
rect 5555 20221 5584 20224
rect 5555 20204 5561 20221
rect 5578 20220 5584 20221
rect 5674 20220 5688 20240
rect 5757 20234 5760 20240
rect 5786 20254 5789 20260
rect 6079 20254 6082 20260
rect 5786 20240 6082 20254
rect 5786 20234 5789 20240
rect 6079 20234 6082 20240
rect 6108 20254 6111 20260
rect 10403 20254 10406 20260
rect 6108 20240 10406 20254
rect 6108 20234 6111 20240
rect 10403 20234 10406 20240
rect 10432 20254 10435 20260
rect 11139 20254 11142 20260
rect 10432 20240 11142 20254
rect 10432 20234 10435 20240
rect 11139 20234 11142 20240
rect 11168 20234 11171 20260
rect 11615 20255 11644 20258
rect 11615 20238 11621 20255
rect 11638 20254 11644 20255
rect 12795 20254 12798 20260
rect 11638 20240 12798 20254
rect 11638 20238 11644 20240
rect 11615 20235 11644 20238
rect 12795 20234 12798 20240
rect 12824 20234 12827 20260
rect 13071 20234 13074 20260
rect 13100 20258 13103 20260
rect 13100 20255 13118 20258
rect 13112 20238 13118 20255
rect 13623 20254 13626 20260
rect 13100 20235 13118 20238
rect 13172 20240 13626 20254
rect 13100 20234 13103 20235
rect 13172 20226 13186 20240
rect 13623 20234 13626 20240
rect 13652 20234 13655 20260
rect 14313 20258 14316 20260
rect 13969 20255 13998 20258
rect 13969 20238 13975 20255
rect 13992 20254 13998 20255
rect 14222 20255 14251 20258
rect 14222 20254 14228 20255
rect 13992 20240 14228 20254
rect 13992 20238 13998 20240
rect 13969 20235 13998 20238
rect 14222 20238 14228 20240
rect 14245 20238 14251 20255
rect 14222 20235 14251 20238
rect 14299 20255 14316 20258
rect 14299 20238 14305 20255
rect 14299 20235 14316 20238
rect 14313 20234 14316 20235
rect 14342 20234 14345 20260
rect 14373 20253 14402 20256
rect 14373 20236 14379 20253
rect 14396 20236 14402 20253
rect 5578 20206 5688 20220
rect 5578 20204 5584 20206
rect 5555 20201 5584 20204
rect 11369 20200 11372 20226
rect 11398 20220 11401 20226
rect 13163 20224 13166 20226
rect 11576 20221 11605 20224
rect 11576 20220 11582 20221
rect 11398 20206 11582 20220
rect 11398 20200 11401 20206
rect 11576 20204 11582 20206
rect 11599 20204 11605 20221
rect 11576 20201 11605 20204
rect 13145 20221 13166 20224
rect 13145 20204 13151 20221
rect 13145 20201 13166 20204
rect 13163 20200 13166 20201
rect 13192 20200 13195 20226
rect 6401 20166 6404 20192
rect 6430 20186 6433 20192
rect 7045 20186 7048 20192
rect 6430 20172 7048 20186
rect 6430 20166 6433 20172
rect 7045 20166 7048 20172
rect 7074 20186 7077 20192
rect 9023 20186 9026 20192
rect 7074 20172 9026 20186
rect 7074 20166 7077 20172
rect 9023 20166 9026 20172
rect 9052 20166 9055 20192
rect 12427 20166 12430 20192
rect 12456 20190 12459 20192
rect 12456 20187 12480 20190
rect 12456 20170 12457 20187
rect 12474 20170 12480 20187
rect 12456 20167 12480 20170
rect 12456 20166 12459 20167
rect 14221 20166 14224 20192
rect 14250 20186 14253 20192
rect 14322 20186 14336 20234
rect 14373 20233 14402 20236
rect 14420 20234 14423 20260
rect 14449 20234 14452 20260
rect 14483 20255 14512 20258
rect 14483 20238 14489 20255
rect 14506 20254 14512 20255
rect 14534 20255 14563 20258
rect 14506 20238 14520 20254
rect 14483 20235 14520 20238
rect 14534 20238 14540 20255
rect 14557 20254 14563 20255
rect 14727 20254 14730 20260
rect 14557 20240 14730 20254
rect 14557 20238 14563 20240
rect 14534 20235 14563 20238
rect 14381 20192 14395 20233
rect 14250 20172 14336 20186
rect 14250 20166 14253 20172
rect 14359 20166 14362 20192
rect 14388 20172 14395 20192
rect 14388 20166 14391 20172
rect 14420 20166 14423 20192
rect 14449 20186 14452 20192
rect 14506 20186 14520 20235
rect 14727 20234 14730 20240
rect 14756 20254 14759 20260
rect 15095 20254 15098 20260
rect 14756 20240 15098 20254
rect 14756 20234 14759 20240
rect 15095 20234 15098 20240
rect 15124 20234 15127 20260
rect 14449 20172 14520 20186
rect 15150 20186 15164 20308
rect 27009 20302 27012 20328
rect 27038 20302 27041 20328
rect 15877 20268 15880 20294
rect 15906 20288 15909 20294
rect 15970 20289 15999 20292
rect 15970 20288 15976 20289
rect 15906 20274 15976 20288
rect 15906 20268 15909 20274
rect 15970 20272 15976 20274
rect 15993 20272 15999 20289
rect 15970 20269 15999 20272
rect 16889 20268 16892 20294
rect 16918 20268 16921 20294
rect 17165 20268 17168 20294
rect 17194 20288 17197 20294
rect 17194 20274 17479 20288
rect 17194 20268 17197 20274
rect 15187 20234 15190 20260
rect 15216 20254 15219 20260
rect 15417 20254 15420 20260
rect 15216 20240 15420 20254
rect 15216 20234 15219 20240
rect 15417 20234 15420 20240
rect 15446 20254 15449 20260
rect 16169 20255 16198 20258
rect 16169 20254 16175 20255
rect 15446 20251 15992 20254
rect 16024 20251 16175 20254
rect 15446 20240 16175 20251
rect 15446 20234 15449 20240
rect 15978 20237 16038 20240
rect 16169 20238 16175 20240
rect 16192 20238 16198 20255
rect 16898 20254 16912 20268
rect 17211 20254 17214 20260
rect 16898 20240 17214 20254
rect 16169 20235 16198 20238
rect 17211 20234 17214 20240
rect 17240 20254 17243 20260
rect 17258 20255 17287 20258
rect 17258 20254 17264 20255
rect 17240 20240 17264 20254
rect 17240 20234 17243 20240
rect 17258 20238 17264 20240
rect 17281 20238 17287 20255
rect 17258 20235 17287 20238
rect 17303 20234 17306 20260
rect 17332 20258 17335 20260
rect 17332 20255 17344 20258
rect 17338 20238 17344 20255
rect 17332 20235 17344 20238
rect 17332 20234 17335 20235
rect 17395 20234 17398 20260
rect 17424 20258 17427 20260
rect 17465 20258 17479 20274
rect 19327 20268 19330 20294
rect 19356 20288 19359 20294
rect 19512 20289 19541 20292
rect 19512 20288 19518 20289
rect 19356 20274 19518 20288
rect 19356 20268 19359 20274
rect 19512 20272 19518 20274
rect 19535 20272 19541 20289
rect 19512 20269 19541 20272
rect 17519 20261 17548 20264
rect 17424 20255 17445 20258
rect 17439 20238 17445 20255
rect 17424 20235 17445 20238
rect 17464 20255 17493 20258
rect 17464 20238 17470 20255
rect 17487 20238 17493 20255
rect 17519 20244 17525 20261
rect 17542 20259 17548 20261
rect 17542 20244 17556 20259
rect 17519 20241 17556 20244
rect 17464 20235 17493 20238
rect 17424 20234 17427 20235
rect 15279 20200 15282 20226
rect 15308 20220 15311 20226
rect 15831 20220 15834 20226
rect 15308 20206 15834 20220
rect 15308 20200 15311 20206
rect 15831 20200 15834 20206
rect 15860 20200 15863 20226
rect 16130 20221 16159 20224
rect 16130 20220 16136 20221
rect 16024 20206 16136 20220
rect 15923 20186 15926 20192
rect 15150 20172 15926 20186
rect 14449 20166 14452 20172
rect 15923 20166 15926 20172
rect 15952 20166 15955 20192
rect 15969 20166 15972 20192
rect 15998 20186 16001 20192
rect 16024 20186 16038 20206
rect 16130 20204 16136 20206
rect 16153 20204 16159 20221
rect 16130 20201 16159 20204
rect 17005 20221 17034 20224
rect 17005 20204 17011 20221
rect 17028 20220 17034 20221
rect 17542 20220 17556 20241
rect 17570 20255 17599 20258
rect 17570 20238 17576 20255
rect 17593 20254 17599 20255
rect 17593 20238 17602 20254
rect 17570 20235 17602 20238
rect 17028 20206 17556 20220
rect 17028 20204 17034 20206
rect 17005 20201 17034 20204
rect 15998 20172 16038 20186
rect 15998 20166 16001 20172
rect 17073 20166 17076 20192
rect 17102 20186 17105 20192
rect 17588 20186 17602 20235
rect 19557 20234 19560 20260
rect 19586 20254 19589 20260
rect 20891 20254 20894 20260
rect 19586 20240 20894 20254
rect 19586 20234 19589 20240
rect 19373 20200 19376 20226
rect 19402 20220 19405 20226
rect 19750 20224 19764 20240
rect 20891 20234 20894 20240
rect 20920 20234 20923 20260
rect 22639 20234 22642 20260
rect 22668 20254 22671 20260
rect 26319 20254 26322 20260
rect 22668 20240 26322 20254
rect 22668 20234 22671 20240
rect 26319 20234 26322 20240
rect 26348 20254 26351 20260
rect 26734 20255 26763 20258
rect 26734 20254 26740 20255
rect 26348 20240 26740 20254
rect 26348 20234 26351 20240
rect 26734 20238 26740 20240
rect 26757 20238 26763 20255
rect 26734 20235 26763 20238
rect 26779 20234 26782 20260
rect 26808 20258 26811 20260
rect 27018 20258 27032 20302
rect 27055 20258 27058 20260
rect 26808 20255 26820 20258
rect 26814 20238 26820 20255
rect 26947 20255 26976 20258
rect 26808 20235 26820 20238
rect 26895 20245 26924 20248
rect 26808 20234 26811 20235
rect 26895 20228 26901 20245
rect 26918 20228 26924 20245
rect 26947 20238 26953 20255
rect 26970 20238 26976 20255
rect 26947 20235 26976 20238
rect 26995 20255 27032 20258
rect 26995 20238 27001 20255
rect 27018 20240 27032 20255
rect 27046 20255 27058 20258
rect 27018 20238 27024 20240
rect 26995 20235 27024 20238
rect 27046 20238 27052 20255
rect 27046 20235 27058 20238
rect 26895 20225 26924 20228
rect 19672 20221 19701 20224
rect 19672 20220 19678 20221
rect 19402 20206 19678 20220
rect 19402 20200 19405 20206
rect 19672 20204 19678 20206
rect 19695 20204 19701 20221
rect 19672 20201 19701 20204
rect 19723 20221 19764 20224
rect 19723 20204 19729 20221
rect 19746 20206 19764 20221
rect 19746 20204 19752 20206
rect 19723 20201 19752 20204
rect 26903 20192 26917 20225
rect 26952 20220 26966 20235
rect 27055 20234 27058 20235
rect 27084 20234 27087 20260
rect 27976 20255 28005 20258
rect 27976 20238 27982 20255
rect 27999 20254 28005 20255
rect 28021 20254 28024 20260
rect 27999 20240 28024 20254
rect 27999 20238 28005 20240
rect 27976 20235 28005 20238
rect 28021 20234 28024 20240
rect 28050 20234 28053 20260
rect 28113 20234 28116 20260
rect 28142 20258 28145 20260
rect 28142 20255 28160 20258
rect 28154 20254 28160 20255
rect 28297 20254 28300 20260
rect 28154 20240 28300 20254
rect 28154 20238 28160 20240
rect 28142 20235 28160 20238
rect 28142 20234 28145 20235
rect 28297 20234 28300 20240
rect 28326 20234 28329 20260
rect 27331 20220 27334 20226
rect 26952 20206 27334 20220
rect 27331 20200 27334 20206
rect 27360 20200 27363 20226
rect 27791 20200 27794 20226
rect 27820 20220 27823 20226
rect 28175 20221 28204 20224
rect 28175 20220 28181 20221
rect 27820 20206 28181 20220
rect 27820 20200 27823 20206
rect 28175 20204 28181 20206
rect 28198 20220 28204 20221
rect 28251 20220 28254 20226
rect 28198 20206 28254 20220
rect 28198 20204 28204 20206
rect 28175 20201 28204 20204
rect 28251 20200 28254 20206
rect 28280 20200 28283 20226
rect 17102 20172 17602 20186
rect 20547 20187 20576 20190
rect 17102 20166 17105 20172
rect 20547 20170 20553 20187
rect 20570 20186 20576 20187
rect 20799 20186 20802 20192
rect 20570 20172 20802 20186
rect 20570 20170 20576 20172
rect 20547 20167 20576 20170
rect 20799 20166 20802 20172
rect 20828 20166 20831 20192
rect 23283 20166 23286 20192
rect 23312 20186 23315 20192
rect 24111 20186 24114 20192
rect 23312 20172 24114 20186
rect 23312 20166 23315 20172
rect 24111 20166 24114 20172
rect 24140 20166 24143 20192
rect 26903 20172 26920 20192
rect 26917 20166 26920 20172
rect 26946 20166 26949 20192
rect 3036 20104 29992 20152
rect 10265 20064 10268 20090
rect 10294 20084 10297 20090
rect 12013 20084 12016 20090
rect 10294 20070 12016 20084
rect 10294 20064 10297 20070
rect 12013 20064 12016 20070
rect 12042 20064 12045 20090
rect 12427 20064 12430 20090
rect 12456 20064 12459 20090
rect 13831 20085 13860 20088
rect 13831 20068 13837 20085
rect 13854 20084 13860 20085
rect 14359 20084 14362 20090
rect 13854 20070 14362 20084
rect 13854 20068 13860 20070
rect 13831 20065 13860 20068
rect 14359 20064 14362 20070
rect 14388 20064 14391 20090
rect 18361 20064 18364 20090
rect 18390 20084 18393 20090
rect 19235 20084 19238 20090
rect 18390 20070 19238 20084
rect 18390 20064 18393 20070
rect 19235 20064 19238 20070
rect 19264 20064 19267 20090
rect 6401 20054 6404 20056
rect 6383 20051 6404 20054
rect 6383 20034 6389 20051
rect 6383 20031 6404 20034
rect 6401 20030 6404 20031
rect 6430 20030 6433 20056
rect 9023 20054 9026 20056
rect 9005 20051 9026 20054
rect 9005 20034 9011 20051
rect 9005 20031 9026 20034
rect 9023 20030 9026 20031
rect 9052 20030 9055 20056
rect 10173 20030 10176 20056
rect 10202 20050 10205 20056
rect 10202 20036 11944 20050
rect 10202 20030 10205 20036
rect 11930 20022 11944 20036
rect 6333 20017 6362 20020
rect 6333 20000 6339 20017
rect 6356 20016 6362 20017
rect 6493 20016 6496 20022
rect 6356 20002 6496 20016
rect 6356 20000 6362 20002
rect 6333 19997 6362 20000
rect 6493 19996 6496 20002
rect 6522 19996 6525 20022
rect 7207 20017 7236 20020
rect 7207 20000 7213 20017
rect 7230 20016 7236 20017
rect 7781 20016 7784 20022
rect 7230 20002 7784 20016
rect 7230 20000 7236 20002
rect 7207 19997 7236 20000
rect 7781 19996 7784 20002
rect 7810 19996 7813 20022
rect 8655 19996 8658 20022
rect 8684 20016 8687 20022
rect 8794 20017 8823 20020
rect 8794 20016 8800 20017
rect 8684 20002 8800 20016
rect 8684 19996 8687 20002
rect 8794 20000 8800 20002
rect 8817 20000 8823 20017
rect 8794 19997 8823 20000
rect 8955 20017 8984 20020
rect 8955 20000 8961 20017
rect 8978 20016 8984 20017
rect 9069 20016 9072 20022
rect 8978 20002 9072 20016
rect 8978 20000 8984 20002
rect 8955 19997 8984 20000
rect 9069 19996 9072 20002
rect 9098 20016 9101 20022
rect 9345 20016 9348 20022
rect 9098 20002 9348 20016
rect 9098 19996 9101 20002
rect 9345 19996 9348 20002
rect 9374 19996 9377 20022
rect 10081 19996 10084 20022
rect 10110 19996 10113 20022
rect 10220 20017 10249 20020
rect 10220 20000 10226 20017
rect 10243 20000 10249 20017
rect 10220 19997 10249 20000
rect 5665 19962 5668 19988
rect 5694 19982 5697 19988
rect 6171 19982 6174 19988
rect 5694 19968 6174 19982
rect 5694 19962 5697 19968
rect 6171 19962 6174 19968
rect 6200 19962 6203 19988
rect 9829 19983 9858 19986
rect 9829 19966 9835 19983
rect 9852 19982 9858 19983
rect 10228 19982 10242 19997
rect 10265 19996 10268 20022
rect 10294 20020 10297 20022
rect 10294 20016 10298 20020
rect 11738 20017 11767 20020
rect 10294 20002 10316 20016
rect 10294 19997 10298 20002
rect 11738 20000 11744 20017
rect 11761 20016 11767 20017
rect 11783 20016 11786 20022
rect 11761 20002 11786 20016
rect 11761 20000 11767 20002
rect 11738 19997 11767 20000
rect 10294 19996 10297 19997
rect 11783 19996 11786 20002
rect 11812 19996 11815 20022
rect 11830 20017 11859 20020
rect 11830 20000 11836 20017
rect 11853 20000 11859 20017
rect 11830 19997 11859 20000
rect 9852 19968 10242 19982
rect 11838 19982 11852 19997
rect 11875 19996 11878 20022
rect 11904 19996 11907 20022
rect 11921 19996 11924 20022
rect 11950 19996 11953 20022
rect 12244 20017 12273 20020
rect 12244 20016 12250 20017
rect 12022 20002 12250 20016
rect 11838 19968 11875 19982
rect 9852 19966 9858 19968
rect 9829 19963 9858 19966
rect 11861 19948 11875 19968
rect 12022 19952 12036 20002
rect 12244 20000 12250 20002
rect 12267 20000 12273 20017
rect 12244 19997 12273 20000
rect 12290 20017 12319 20020
rect 12290 20000 12296 20017
rect 12313 20016 12319 20017
rect 12335 20016 12338 20022
rect 12313 20002 12338 20016
rect 12313 20000 12319 20002
rect 12290 19997 12319 20000
rect 12335 19996 12338 20002
rect 12364 19996 12367 20022
rect 12381 19996 12384 20022
rect 12410 19996 12413 20022
rect 12436 20020 12450 20064
rect 12611 20030 12614 20056
rect 12640 20050 12643 20056
rect 13025 20054 13028 20056
rect 12956 20051 12985 20054
rect 12956 20050 12962 20051
rect 12640 20036 12962 20050
rect 12640 20030 12643 20036
rect 12956 20034 12962 20036
rect 12979 20034 12985 20051
rect 12956 20031 12985 20034
rect 13007 20051 13028 20054
rect 13007 20034 13013 20051
rect 13007 20031 13028 20034
rect 13025 20030 13028 20031
rect 13054 20030 13057 20056
rect 15601 20030 15604 20056
rect 15630 20050 15633 20056
rect 15763 20051 15792 20054
rect 15763 20050 15769 20051
rect 15630 20036 15769 20050
rect 15630 20030 15633 20036
rect 15763 20034 15769 20036
rect 15786 20034 15792 20051
rect 15763 20031 15792 20034
rect 17929 20051 17958 20054
rect 17929 20034 17935 20051
rect 17952 20050 17958 20051
rect 17952 20036 18062 20050
rect 17952 20034 17958 20036
rect 17929 20031 17958 20034
rect 12428 20017 12457 20020
rect 12428 20000 12434 20017
rect 12451 20000 12457 20017
rect 12428 19997 12457 20000
rect 12488 20017 12517 20020
rect 12488 20000 12494 20017
rect 12511 20016 12517 20017
rect 12511 20002 12634 20016
rect 12511 20000 12517 20002
rect 12488 19997 12517 20000
rect 12620 19988 12634 20002
rect 13117 19996 13120 20022
rect 13146 20016 13149 20022
rect 15003 20016 15006 20022
rect 13146 20002 15006 20016
rect 13146 19996 13149 20002
rect 15003 19996 15006 20002
rect 15032 19996 15035 20022
rect 15141 19996 15144 20022
rect 15170 20016 15173 20022
rect 15711 20017 15740 20020
rect 15711 20016 15717 20017
rect 15170 20002 15717 20016
rect 15170 19996 15173 20002
rect 15711 20000 15717 20002
rect 15734 20016 15740 20017
rect 15969 20016 15972 20022
rect 15734 20002 15972 20016
rect 15734 20000 15740 20002
rect 15711 19997 15740 20000
rect 15969 19996 15972 20002
rect 15998 20016 16001 20022
rect 16107 20016 16110 20022
rect 15998 20002 16110 20016
rect 15998 19996 16001 20002
rect 16107 19996 16110 20002
rect 16136 19996 16139 20022
rect 16591 20017 16620 20020
rect 16591 20000 16597 20017
rect 16614 20016 16620 20017
rect 17303 20016 17306 20022
rect 16614 20002 17306 20016
rect 16614 20000 16620 20002
rect 16591 19997 16620 20000
rect 17303 19996 17306 20002
rect 17332 19996 17335 20022
rect 17855 19996 17858 20022
rect 17884 20020 17887 20022
rect 17884 20017 17902 20020
rect 17896 20000 17902 20017
rect 18048 20016 18062 20036
rect 19060 20036 19166 20050
rect 18361 20016 18364 20022
rect 18048 20002 18364 20016
rect 17884 19997 17902 20000
rect 17884 19996 17887 19997
rect 18361 19996 18364 20002
rect 18390 19996 18393 20022
rect 19006 20017 19035 20020
rect 19006 20000 19012 20017
rect 19029 20016 19035 20017
rect 19060 20016 19074 20036
rect 19029 20002 19074 20016
rect 19098 20017 19127 20020
rect 19029 20000 19035 20002
rect 19006 19997 19035 20000
rect 19098 20000 19104 20017
rect 19121 20000 19127 20017
rect 19152 20016 19166 20036
rect 20799 20030 20802 20056
rect 20828 20030 20831 20056
rect 23219 20051 23248 20054
rect 23219 20034 23225 20051
rect 23242 20050 23248 20051
rect 23283 20050 23286 20056
rect 23242 20036 23286 20050
rect 23242 20034 23248 20036
rect 23219 20031 23248 20034
rect 23283 20030 23286 20036
rect 23312 20030 23315 20056
rect 24111 20030 24114 20056
rect 24140 20050 24143 20056
rect 25783 20051 25812 20054
rect 25783 20050 25789 20051
rect 24140 20036 25789 20050
rect 24140 20030 24143 20036
rect 25783 20034 25789 20036
rect 25806 20034 25812 20051
rect 25783 20031 25812 20034
rect 20339 20016 20342 20022
rect 19152 20002 20342 20016
rect 19098 19997 19127 20000
rect 12611 19962 12614 19988
rect 12640 19962 12643 19988
rect 12749 19962 12752 19988
rect 12778 19982 12781 19988
rect 12796 19983 12825 19986
rect 12796 19982 12802 19983
rect 12778 19968 12802 19982
rect 12778 19962 12781 19968
rect 12796 19966 12802 19968
rect 12819 19966 12825 19983
rect 12796 19963 12825 19966
rect 15556 19983 15585 19986
rect 15556 19966 15562 19983
rect 15579 19966 15585 19983
rect 15556 19963 15585 19966
rect 9653 19934 11875 19948
rect 9345 19894 9348 19920
rect 9374 19914 9377 19920
rect 9653 19914 9667 19934
rect 9374 19900 9667 19914
rect 10082 19915 10111 19918
rect 9374 19894 9377 19900
rect 10082 19898 10088 19915
rect 10105 19914 10111 19915
rect 10311 19914 10314 19920
rect 10105 19900 10314 19914
rect 10105 19898 10111 19900
rect 10082 19895 10111 19898
rect 10311 19894 10314 19900
rect 10340 19894 10343 19920
rect 11861 19914 11875 19934
rect 12014 19949 12043 19952
rect 12014 19932 12020 19949
rect 12037 19932 12043 19949
rect 12014 19929 12043 19932
rect 12244 19949 12273 19952
rect 12244 19932 12250 19949
rect 12267 19948 12273 19949
rect 12703 19948 12706 19954
rect 12267 19934 12706 19948
rect 12267 19932 12273 19934
rect 12244 19929 12273 19932
rect 12703 19928 12706 19934
rect 12732 19928 12735 19954
rect 12059 19914 12062 19920
rect 11861 19900 12062 19914
rect 12059 19894 12062 19900
rect 12088 19894 12091 19920
rect 15564 19914 15578 19963
rect 17717 19962 17720 19988
rect 17746 19962 17749 19988
rect 18753 19983 18782 19986
rect 18753 19966 18759 19983
rect 18776 19982 18782 19983
rect 19106 19982 19120 19997
rect 20339 19996 20342 20002
rect 20368 19996 20371 20022
rect 20569 19996 20572 20022
rect 20598 20016 20601 20022
rect 20616 20017 20645 20020
rect 20616 20016 20622 20017
rect 20598 20002 20622 20016
rect 20598 19996 20601 20002
rect 20616 20000 20622 20002
rect 20639 20000 20645 20017
rect 20616 19997 20645 20000
rect 20661 19996 20664 20022
rect 20690 19996 20693 20022
rect 20753 19996 20756 20022
rect 20782 19996 20785 20022
rect 20846 20017 20875 20020
rect 20846 20000 20852 20017
rect 20869 20016 20875 20017
rect 20937 20016 20940 20022
rect 20869 20002 20940 20016
rect 20869 20000 20875 20002
rect 20846 19997 20875 20000
rect 20937 19996 20940 20002
rect 20966 20016 20969 20022
rect 22685 20016 22688 20022
rect 20966 20002 22688 20016
rect 20966 19996 20969 20002
rect 22685 19996 22688 20002
rect 22714 19996 22717 20022
rect 23008 20017 23037 20020
rect 23008 20000 23014 20017
rect 23031 20016 23037 20017
rect 23053 20016 23056 20022
rect 23031 20002 23056 20016
rect 23031 20000 23037 20002
rect 23008 19997 23037 20000
rect 23053 19996 23056 20002
rect 23082 19996 23085 20022
rect 23145 19996 23148 20022
rect 23174 20020 23177 20022
rect 23174 20017 23192 20020
rect 23186 20016 23192 20017
rect 23559 20016 23562 20022
rect 23186 20002 23562 20016
rect 23186 20000 23192 20002
rect 23174 19997 23192 20000
rect 23174 19996 23177 19997
rect 23559 19996 23562 20002
rect 23588 19996 23591 20022
rect 24043 20017 24072 20020
rect 24043 20000 24049 20017
rect 24066 20016 24072 20017
rect 24296 20017 24325 20020
rect 24296 20016 24302 20017
rect 24066 20002 24302 20016
rect 24066 20000 24072 20002
rect 24043 19997 24072 20000
rect 24296 20000 24302 20002
rect 24319 20000 24325 20017
rect 24388 20017 24417 20020
rect 24388 20016 24394 20017
rect 24296 19997 24325 20000
rect 24350 20002 24394 20016
rect 24350 19982 24364 20002
rect 24388 20000 24394 20002
rect 24411 20000 24417 20017
rect 24388 19997 24417 20000
rect 24433 19996 24436 20022
rect 24462 19996 24465 20022
rect 24479 19996 24482 20022
rect 24508 20020 24511 20022
rect 24508 20016 24512 20020
rect 24508 20002 24530 20016
rect 24508 19997 24512 20002
rect 24508 19996 24511 19997
rect 25537 19996 25540 20022
rect 25566 20016 25569 20022
rect 25584 20017 25613 20020
rect 25584 20016 25590 20017
rect 25566 20002 25590 20016
rect 25566 19996 25569 20002
rect 25584 20000 25590 20002
rect 25607 20000 25613 20017
rect 25584 19997 25613 20000
rect 25721 19996 25724 20022
rect 25750 20020 25753 20022
rect 25750 20017 25768 20020
rect 25762 20000 25768 20017
rect 25750 19997 25768 20000
rect 26619 20017 26648 20020
rect 26619 20000 26625 20017
rect 26642 20016 26648 20017
rect 26917 20016 26920 20022
rect 26642 20002 26920 20016
rect 26642 20000 26648 20002
rect 26619 19997 26648 20000
rect 25750 19996 25753 19997
rect 26917 19996 26920 20002
rect 26946 19996 26949 20022
rect 18776 19968 19120 19982
rect 24258 19968 24364 19982
rect 18776 19966 18782 19968
rect 18753 19963 18782 19966
rect 20891 19928 20894 19954
rect 20920 19948 20923 19954
rect 22961 19948 22964 19954
rect 20920 19934 22964 19948
rect 20920 19928 20923 19934
rect 22961 19928 22964 19934
rect 22990 19928 22993 19954
rect 24258 19920 24272 19968
rect 15877 19914 15880 19920
rect 15564 19900 15880 19914
rect 15877 19894 15880 19900
rect 15906 19914 15909 19920
rect 15969 19914 15972 19920
rect 15906 19900 15972 19914
rect 15906 19894 15909 19900
rect 15969 19894 15972 19900
rect 15998 19894 16001 19920
rect 18867 19894 18870 19920
rect 18896 19914 18899 19920
rect 19052 19915 19081 19918
rect 19052 19914 19058 19915
rect 18896 19900 19058 19914
rect 18896 19894 18899 19900
rect 19052 19898 19058 19900
rect 19075 19898 19081 19915
rect 19052 19895 19081 19898
rect 20616 19915 20645 19918
rect 20616 19898 20622 19915
rect 20639 19914 20645 19915
rect 20661 19914 20664 19920
rect 20639 19900 20664 19914
rect 20639 19898 20645 19900
rect 20616 19895 20645 19898
rect 20661 19894 20664 19900
rect 20690 19894 20693 19920
rect 23099 19894 23102 19920
rect 23128 19914 23131 19920
rect 24249 19914 24252 19920
rect 23128 19900 24252 19914
rect 23128 19894 23131 19900
rect 24249 19894 24252 19900
rect 24278 19894 24281 19920
rect 24295 19894 24298 19920
rect 24324 19894 24327 19920
rect 24479 19894 24482 19920
rect 24508 19914 24511 19920
rect 29263 19914 29266 19920
rect 24508 19900 29266 19914
rect 24508 19894 24511 19900
rect 29263 19894 29266 19900
rect 29292 19894 29295 19920
rect 3036 19832 29992 19880
rect 5665 19812 5668 19818
rect 5398 19798 5668 19812
rect 5343 19724 5346 19750
rect 5372 19744 5375 19750
rect 5398 19748 5412 19798
rect 5665 19792 5668 19798
rect 5694 19792 5697 19818
rect 9691 19813 9720 19816
rect 9691 19796 9697 19813
rect 9714 19812 9720 19813
rect 10081 19812 10084 19818
rect 9714 19798 10084 19812
rect 9714 19796 9720 19798
rect 9691 19793 9720 19796
rect 10081 19792 10084 19798
rect 10110 19792 10113 19818
rect 11047 19812 11050 19818
rect 10964 19798 11050 19812
rect 5390 19745 5419 19748
rect 5390 19744 5396 19745
rect 5372 19730 5396 19744
rect 5372 19724 5375 19730
rect 5390 19728 5396 19730
rect 5413 19728 5419 19745
rect 5390 19725 5419 19728
rect 8655 19724 8658 19750
rect 8684 19724 8687 19750
rect 9575 19724 9578 19750
rect 9604 19744 9607 19750
rect 10220 19745 10249 19748
rect 10220 19744 10226 19745
rect 9604 19730 10226 19744
rect 9604 19724 9607 19730
rect 10220 19728 10226 19730
rect 10243 19728 10249 19745
rect 10220 19725 10249 19728
rect 10588 19745 10617 19748
rect 10588 19728 10594 19745
rect 10611 19744 10617 19745
rect 10725 19744 10728 19750
rect 10611 19730 10728 19744
rect 10611 19728 10617 19730
rect 10588 19725 10617 19728
rect 10725 19724 10728 19730
rect 10754 19724 10757 19750
rect 10964 19748 10978 19798
rect 11047 19792 11050 19798
rect 11076 19792 11079 19818
rect 11875 19792 11878 19818
rect 11904 19812 11907 19818
rect 11991 19813 12020 19816
rect 11991 19812 11997 19813
rect 11904 19798 11997 19812
rect 11904 19792 11907 19798
rect 11991 19796 11997 19798
rect 12014 19796 12020 19813
rect 11991 19793 12020 19796
rect 12059 19792 12062 19818
rect 12088 19812 12091 19818
rect 14015 19813 14044 19816
rect 12088 19798 13830 19812
rect 12088 19792 12091 19798
rect 12519 19758 12522 19784
rect 12548 19778 12551 19784
rect 12611 19778 12614 19784
rect 12548 19764 12614 19778
rect 12548 19758 12551 19764
rect 12611 19758 12614 19764
rect 12640 19758 12643 19784
rect 13816 19778 13830 19798
rect 14015 19796 14021 19813
rect 14038 19812 14044 19813
rect 14359 19812 14362 19818
rect 14038 19798 14362 19812
rect 14038 19796 14044 19798
rect 14015 19793 14044 19796
rect 14359 19792 14362 19798
rect 14388 19792 14391 19818
rect 17005 19813 17034 19816
rect 17005 19796 17011 19813
rect 17028 19812 17034 19813
rect 17395 19812 17398 19818
rect 17028 19798 17398 19812
rect 17028 19796 17034 19798
rect 17005 19793 17034 19796
rect 17395 19792 17398 19798
rect 17424 19792 17427 19818
rect 21443 19812 21446 19818
rect 20693 19798 21446 19812
rect 14727 19778 14730 19784
rect 13816 19764 14730 19778
rect 14727 19758 14730 19764
rect 14756 19758 14759 19784
rect 10956 19745 10985 19748
rect 10956 19728 10962 19745
rect 10979 19728 10985 19745
rect 10956 19725 10985 19728
rect 19327 19724 19330 19750
rect 19356 19744 19359 19750
rect 19374 19745 19403 19748
rect 19374 19744 19380 19745
rect 19356 19730 19380 19744
rect 19356 19724 19359 19730
rect 19374 19728 19380 19730
rect 19397 19728 19403 19745
rect 19374 19725 19403 19728
rect 5527 19690 5530 19716
rect 5556 19714 5559 19716
rect 5556 19711 5574 19714
rect 5568 19694 5574 19711
rect 5556 19691 5574 19694
rect 8817 19711 8846 19714
rect 8817 19694 8823 19711
rect 8840 19710 8846 19711
rect 9069 19710 9072 19716
rect 8840 19696 9072 19710
rect 8840 19694 8846 19696
rect 8817 19691 8846 19694
rect 5556 19690 5559 19691
rect 9069 19690 9072 19696
rect 9098 19690 9101 19716
rect 10311 19690 10314 19716
rect 10340 19690 10343 19716
rect 10357 19690 10360 19716
rect 10386 19690 10389 19716
rect 11117 19711 11146 19714
rect 11117 19694 11123 19711
rect 11140 19710 11146 19711
rect 11369 19710 11372 19716
rect 11140 19696 11372 19710
rect 11140 19694 11146 19696
rect 11117 19691 11146 19694
rect 11369 19690 11372 19696
rect 11398 19690 11401 19716
rect 12749 19690 12752 19716
rect 12778 19710 12781 19716
rect 12980 19711 13009 19714
rect 12980 19710 12986 19711
rect 12778 19696 12986 19710
rect 12778 19690 12781 19696
rect 12980 19694 12986 19696
rect 13003 19694 13009 19711
rect 12980 19691 13009 19694
rect 13025 19690 13028 19716
rect 13054 19710 13057 19716
rect 13179 19711 13208 19714
rect 13179 19710 13185 19711
rect 13054 19696 13185 19710
rect 13054 19690 13057 19696
rect 13179 19694 13185 19696
rect 13202 19710 13208 19711
rect 13301 19710 13304 19716
rect 13202 19696 13304 19710
rect 13202 19694 13208 19696
rect 13179 19691 13208 19694
rect 13301 19690 13304 19696
rect 13330 19690 13333 19716
rect 15969 19690 15972 19716
rect 15998 19690 16001 19716
rect 16107 19690 16110 19716
rect 16136 19714 16139 19716
rect 16136 19711 16154 19714
rect 16148 19694 16154 19711
rect 20693 19710 20707 19798
rect 21443 19792 21446 19798
rect 21472 19792 21475 19818
rect 24249 19792 24252 19818
rect 24278 19812 24281 19818
rect 27331 19812 27334 19818
rect 24278 19798 27334 19812
rect 24278 19792 24281 19798
rect 27331 19792 27334 19798
rect 27360 19792 27363 19818
rect 22685 19758 22688 19784
rect 22714 19778 22717 19784
rect 24479 19778 24482 19784
rect 22714 19764 24482 19778
rect 22714 19758 22717 19764
rect 24479 19758 24482 19764
rect 24508 19758 24511 19784
rect 16136 19691 16154 19694
rect 19704 19696 20707 19710
rect 16136 19690 16139 19691
rect 5619 19680 5622 19682
rect 5601 19677 5622 19680
rect 5601 19660 5607 19677
rect 5601 19657 5622 19660
rect 5619 19656 5622 19657
rect 5648 19656 5651 19682
rect 8701 19656 8704 19682
rect 8730 19676 8733 19682
rect 11185 19680 11188 19682
rect 8863 19677 8892 19680
rect 8863 19676 8869 19677
rect 8730 19662 8869 19676
rect 8730 19656 8733 19662
rect 8863 19660 8869 19662
rect 8886 19660 8892 19677
rect 8863 19657 8892 19660
rect 11167 19677 11188 19680
rect 11167 19660 11173 19677
rect 11167 19657 11188 19660
rect 11185 19656 11188 19657
rect 11214 19656 11217 19682
rect 13140 19677 13169 19680
rect 13140 19676 13146 19677
rect 12988 19662 13146 19676
rect 12988 19648 13002 19662
rect 13140 19660 13146 19662
rect 13163 19660 13169 19677
rect 13140 19657 13169 19660
rect 16181 19677 16210 19680
rect 16181 19660 16187 19677
rect 16204 19676 16210 19677
rect 16245 19676 16248 19682
rect 16204 19662 16248 19676
rect 16204 19660 16210 19662
rect 16181 19657 16210 19660
rect 16245 19656 16248 19662
rect 16274 19656 16277 19682
rect 19373 19656 19376 19682
rect 19402 19676 19405 19682
rect 19534 19677 19563 19680
rect 19534 19676 19540 19677
rect 19402 19662 19540 19676
rect 19402 19656 19405 19662
rect 19534 19660 19540 19662
rect 19557 19660 19563 19677
rect 19534 19657 19563 19660
rect 19585 19677 19614 19680
rect 19585 19660 19591 19677
rect 19608 19676 19614 19677
rect 19704 19676 19718 19696
rect 21075 19690 21078 19716
rect 21104 19710 21107 19716
rect 21259 19710 21262 19716
rect 21104 19696 21262 19710
rect 21104 19690 21107 19696
rect 21259 19690 21262 19696
rect 21288 19710 21291 19716
rect 21306 19711 21335 19714
rect 21306 19710 21312 19711
rect 21288 19696 21312 19710
rect 21288 19690 21291 19696
rect 21306 19694 21312 19696
rect 21329 19694 21335 19711
rect 21306 19691 21335 19694
rect 21505 19711 21534 19714
rect 21505 19694 21511 19711
rect 21528 19710 21534 19711
rect 21581 19710 21584 19716
rect 21528 19696 21584 19710
rect 21528 19694 21534 19696
rect 21505 19691 21534 19694
rect 21581 19690 21584 19696
rect 21610 19710 21613 19716
rect 23283 19710 23286 19716
rect 21610 19696 23286 19710
rect 21610 19690 21613 19696
rect 23283 19690 23286 19696
rect 23312 19690 23315 19716
rect 19608 19662 19718 19676
rect 19608 19660 19614 19662
rect 19585 19657 19614 19660
rect 21351 19656 21354 19682
rect 21380 19676 21383 19682
rect 21466 19677 21495 19680
rect 21466 19676 21472 19677
rect 21380 19662 21472 19676
rect 21380 19656 21383 19662
rect 21466 19660 21472 19662
rect 21489 19660 21495 19677
rect 21466 19657 21495 19660
rect 6401 19622 6404 19648
rect 6430 19646 6433 19648
rect 6430 19643 6454 19646
rect 6430 19626 6431 19643
rect 6448 19626 6454 19643
rect 6430 19623 6454 19626
rect 6430 19622 6433 19623
rect 12979 19622 12982 19648
rect 13008 19622 13011 19648
rect 20431 19646 20434 19648
rect 20409 19643 20434 19646
rect 20409 19626 20415 19643
rect 20432 19626 20434 19643
rect 20409 19623 20434 19626
rect 20431 19622 20434 19623
rect 20460 19622 20463 19648
rect 22341 19643 22370 19646
rect 22341 19626 22347 19643
rect 22364 19642 22370 19643
rect 22731 19642 22734 19648
rect 22364 19628 22734 19642
rect 22364 19626 22370 19628
rect 22341 19623 22370 19626
rect 22731 19622 22734 19628
rect 22760 19622 22763 19648
rect 22961 19622 22964 19648
rect 22990 19642 22993 19648
rect 27791 19642 27794 19648
rect 22990 19628 27794 19642
rect 22990 19622 22993 19628
rect 27791 19622 27794 19628
rect 27820 19622 27823 19648
rect 3036 19560 29992 19608
rect 11185 19520 11188 19546
rect 11214 19540 11217 19546
rect 12611 19540 12614 19546
rect 11214 19526 12614 19540
rect 11214 19520 11217 19526
rect 12611 19520 12614 19526
rect 12640 19540 12643 19546
rect 13163 19540 13166 19546
rect 12640 19526 13166 19540
rect 12640 19520 12643 19526
rect 13163 19520 13166 19526
rect 13192 19520 13195 19546
rect 20569 19520 20572 19546
rect 20598 19520 20601 19546
rect 22593 19520 22596 19546
rect 22622 19520 22625 19546
rect 22777 19520 22780 19546
rect 22806 19540 22809 19546
rect 24181 19541 24210 19544
rect 22806 19526 22869 19540
rect 22806 19520 22809 19526
rect 3779 19510 3782 19512
rect 3761 19507 3782 19510
rect 3761 19490 3767 19507
rect 3761 19487 3782 19490
rect 3779 19486 3782 19487
rect 3808 19486 3811 19512
rect 4975 19486 4978 19512
rect 5004 19506 5007 19512
rect 7487 19507 7516 19510
rect 5004 19487 5016 19506
rect 7487 19490 7493 19507
rect 7510 19506 7516 19507
rect 7551 19506 7554 19512
rect 7510 19492 7554 19506
rect 7510 19490 7516 19492
rect 7487 19487 7516 19490
rect 5004 19486 5028 19487
rect 4999 19484 5028 19486
rect 3549 19452 3552 19478
rect 3578 19452 3581 19478
rect 3595 19452 3598 19478
rect 3624 19472 3627 19478
rect 3711 19473 3740 19476
rect 3711 19472 3717 19473
rect 3624 19458 3717 19472
rect 3624 19452 3627 19458
rect 3711 19456 3717 19458
rect 3734 19472 3740 19473
rect 3734 19458 4538 19472
rect 3734 19456 3740 19458
rect 3711 19453 3740 19456
rect 4524 19404 4538 19458
rect 4837 19452 4840 19478
rect 4866 19452 4869 19478
rect 4929 19476 4932 19478
rect 4915 19473 4932 19476
rect 4915 19456 4921 19473
rect 4915 19453 4932 19456
rect 4929 19452 4932 19453
rect 4958 19452 4961 19478
rect 4999 19467 5005 19484
rect 5022 19467 5028 19484
rect 4999 19464 5028 19467
rect 5044 19484 5073 19487
rect 7551 19486 7554 19492
rect 7580 19486 7583 19512
rect 8311 19507 8340 19510
rect 8311 19490 8317 19507
rect 8334 19506 8340 19507
rect 8334 19492 9077 19506
rect 8334 19490 8340 19492
rect 8311 19487 8340 19490
rect 5044 19467 5050 19484
rect 5067 19467 5073 19484
rect 5159 19476 5162 19478
rect 5044 19464 5073 19467
rect 5099 19473 5128 19476
rect 5045 19444 5059 19464
rect 5099 19456 5105 19473
rect 5122 19456 5128 19473
rect 5099 19453 5128 19456
rect 5150 19473 5162 19476
rect 5150 19456 5156 19473
rect 5150 19453 5162 19456
rect 4585 19439 4614 19442
rect 4585 19422 4591 19439
rect 4608 19438 4614 19439
rect 4608 19424 4998 19438
rect 4608 19422 4614 19424
rect 4585 19419 4614 19422
rect 4929 19404 4932 19410
rect 4524 19390 4932 19404
rect 4929 19384 4932 19390
rect 4958 19384 4961 19410
rect 4984 19404 4998 19424
rect 5021 19418 5024 19444
rect 5050 19424 5059 19444
rect 5050 19418 5053 19424
rect 4984 19390 5059 19404
rect 4837 19350 4840 19376
rect 4866 19350 4869 19376
rect 5045 19370 5059 19390
rect 5107 19370 5121 19453
rect 5159 19452 5162 19453
rect 5188 19452 5191 19478
rect 7275 19452 7278 19478
rect 7304 19452 7307 19478
rect 7413 19452 7416 19478
rect 7442 19476 7445 19478
rect 7442 19473 7460 19476
rect 7454 19456 7460 19473
rect 7442 19453 7460 19456
rect 7442 19452 7445 19453
rect 8379 19452 8382 19478
rect 8408 19472 8411 19478
rect 8794 19473 8823 19476
rect 8794 19472 8800 19473
rect 8408 19458 8800 19472
rect 8408 19452 8411 19458
rect 8794 19456 8800 19458
rect 8817 19456 8823 19473
rect 8794 19453 8823 19456
rect 8802 19438 8816 19453
rect 8839 19452 8842 19478
rect 8868 19476 8871 19478
rect 9063 19476 9077 19492
rect 20063 19486 20066 19512
rect 20092 19506 20095 19512
rect 20386 19507 20415 19510
rect 20386 19506 20392 19507
rect 20092 19492 20392 19506
rect 20092 19486 20095 19492
rect 20386 19490 20392 19492
rect 20409 19490 20415 19507
rect 20386 19487 20415 19490
rect 20431 19486 20434 19512
rect 20460 19486 20463 19512
rect 21305 19510 21308 19512
rect 21287 19507 21308 19510
rect 21287 19490 21293 19507
rect 21287 19487 21308 19490
rect 21305 19486 21308 19487
rect 21334 19486 21337 19512
rect 22855 19487 22869 19526
rect 24181 19524 24187 19541
rect 24204 19540 24210 19541
rect 24433 19540 24436 19546
rect 24204 19526 24436 19540
rect 24204 19524 24210 19526
rect 24181 19521 24210 19524
rect 24433 19520 24436 19526
rect 24462 19520 24465 19546
rect 22847 19484 22876 19487
rect 22961 19486 22964 19512
rect 22990 19506 22993 19512
rect 23345 19507 23374 19510
rect 23345 19506 23351 19507
rect 22990 19492 23351 19506
rect 22990 19486 22993 19492
rect 23345 19490 23351 19492
rect 23368 19490 23374 19507
rect 23345 19487 23374 19490
rect 9115 19476 9118 19478
rect 8868 19473 8880 19476
rect 8874 19456 8880 19473
rect 9007 19473 9036 19476
rect 8868 19453 8880 19456
rect 8955 19468 8984 19471
rect 8868 19452 8871 19453
rect 8955 19451 8961 19468
rect 8978 19451 8984 19468
rect 9007 19456 9013 19473
rect 9030 19456 9036 19473
rect 9007 19453 9036 19456
rect 9055 19473 9084 19476
rect 9055 19456 9061 19473
rect 9078 19456 9084 19473
rect 9055 19453 9084 19456
rect 9106 19473 9118 19476
rect 9106 19456 9112 19473
rect 9144 19472 9147 19478
rect 9207 19472 9210 19478
rect 9144 19458 9210 19472
rect 9106 19453 9118 19456
rect 8955 19448 8984 19451
rect 8802 19424 8862 19438
rect 8241 19384 8244 19410
rect 8270 19404 8273 19410
rect 8794 19405 8823 19408
rect 8794 19404 8800 19405
rect 8270 19390 8800 19404
rect 8270 19384 8273 19390
rect 8794 19388 8800 19390
rect 8817 19388 8823 19405
rect 8794 19385 8823 19388
rect 5045 19356 5121 19370
rect 8848 19370 8862 19424
rect 8963 19410 8977 19448
rect 9015 19438 9029 19453
rect 9115 19452 9118 19453
rect 9144 19452 9147 19458
rect 9207 19452 9210 19458
rect 9236 19472 9239 19478
rect 12519 19472 12522 19478
rect 9236 19458 12522 19472
rect 9236 19452 9239 19458
rect 12519 19452 12522 19458
rect 12548 19452 12551 19478
rect 20293 19452 20296 19478
rect 20322 19452 20325 19478
rect 20478 19473 20507 19476
rect 20478 19456 20484 19473
rect 20501 19472 20507 19473
rect 20501 19458 20707 19472
rect 20501 19456 20507 19458
rect 20478 19453 20507 19456
rect 9299 19438 9302 19444
rect 9015 19424 9302 19438
rect 9299 19418 9302 19424
rect 9328 19438 9331 19444
rect 9621 19438 9624 19444
rect 9328 19424 9624 19438
rect 9328 19418 9331 19424
rect 9621 19418 9624 19424
rect 9650 19418 9653 19444
rect 8963 19390 8980 19410
rect 8977 19384 8980 19390
rect 9006 19384 9009 19410
rect 9299 19370 9302 19376
rect 8848 19356 9302 19370
rect 9299 19350 9302 19356
rect 9328 19370 9331 19376
rect 12381 19370 12384 19376
rect 9328 19356 12384 19370
rect 9328 19350 9331 19356
rect 12381 19350 12384 19356
rect 12410 19350 12413 19376
rect 20693 19370 20707 19458
rect 21029 19452 21032 19478
rect 21058 19472 21061 19478
rect 21231 19473 21260 19476
rect 21231 19472 21237 19473
rect 21058 19458 21237 19472
rect 21058 19452 21061 19458
rect 21231 19456 21237 19458
rect 21254 19472 21260 19473
rect 21351 19472 21354 19478
rect 21254 19458 21354 19472
rect 21254 19456 21260 19458
rect 21231 19453 21260 19456
rect 21351 19452 21354 19458
rect 21380 19452 21383 19478
rect 22593 19452 22596 19478
rect 22622 19452 22625 19478
rect 22651 19473 22680 19476
rect 22651 19472 22657 19473
rect 22648 19456 22657 19472
rect 22674 19456 22680 19473
rect 22648 19453 22680 19456
rect 21075 19418 21078 19444
rect 21104 19418 21107 19444
rect 22111 19439 22140 19442
rect 22111 19422 22117 19439
rect 22134 19438 22140 19439
rect 22648 19438 22662 19453
rect 22731 19452 22734 19478
rect 22760 19476 22763 19478
rect 22760 19473 22774 19476
rect 22768 19456 22774 19473
rect 22760 19453 22774 19456
rect 22793 19473 22822 19476
rect 22793 19456 22799 19473
rect 22816 19456 22822 19473
rect 22847 19467 22853 19484
rect 22870 19467 22876 19484
rect 22915 19476 22918 19478
rect 22847 19464 22876 19467
rect 22906 19473 22918 19476
rect 22793 19453 22822 19456
rect 22906 19456 22912 19473
rect 22906 19453 22918 19456
rect 22760 19452 22763 19453
rect 22134 19424 22662 19438
rect 22801 19438 22815 19453
rect 22915 19452 22918 19453
rect 22944 19452 22947 19478
rect 23191 19452 23194 19478
rect 23220 19472 23223 19478
rect 23301 19473 23330 19476
rect 23301 19472 23307 19473
rect 23220 19458 23307 19472
rect 23220 19452 23223 19458
rect 23301 19456 23307 19458
rect 23324 19456 23330 19473
rect 23301 19453 23330 19456
rect 22801 19424 22846 19438
rect 22134 19422 22140 19424
rect 22111 19419 22140 19422
rect 22832 19376 22846 19424
rect 22961 19418 22964 19444
rect 22990 19438 22993 19444
rect 23053 19438 23056 19444
rect 22990 19424 23056 19438
rect 22990 19418 22993 19424
rect 23053 19418 23056 19424
rect 23082 19438 23085 19444
rect 23146 19439 23175 19442
rect 23146 19438 23152 19439
rect 23082 19424 23152 19438
rect 23082 19418 23085 19424
rect 23146 19422 23152 19424
rect 23169 19422 23175 19439
rect 23146 19419 23175 19422
rect 22639 19370 22642 19376
rect 20693 19356 22642 19370
rect 22639 19350 22642 19356
rect 22668 19350 22671 19376
rect 22823 19350 22826 19376
rect 22852 19370 22855 19376
rect 23099 19370 23102 19376
rect 22852 19356 23102 19370
rect 22852 19350 22855 19356
rect 23099 19350 23102 19356
rect 23128 19350 23131 19376
rect 3036 19288 29992 19336
rect 4171 19269 4200 19272
rect 4171 19252 4177 19269
rect 4194 19268 4200 19269
rect 4883 19268 4886 19274
rect 4194 19254 4886 19268
rect 4194 19252 4200 19254
rect 4171 19249 4200 19252
rect 4883 19248 4886 19254
rect 4912 19248 4915 19274
rect 5665 19268 5668 19274
rect 5536 19254 5668 19268
rect 5536 19204 5550 19254
rect 5665 19248 5668 19254
rect 5694 19248 5697 19274
rect 5803 19248 5806 19274
rect 5832 19268 5835 19274
rect 6862 19269 6891 19272
rect 6862 19268 6868 19269
rect 5832 19254 6868 19268
rect 5832 19248 5835 19254
rect 6862 19252 6868 19254
rect 6885 19252 6891 19269
rect 8241 19268 8244 19274
rect 6862 19249 6891 19252
rect 6962 19254 8244 19268
rect 5528 19201 5557 19204
rect 5528 19184 5534 19201
rect 5551 19184 5557 19201
rect 5528 19181 5557 19184
rect 3135 19146 3138 19172
rect 3164 19146 3167 19172
rect 3297 19167 3326 19170
rect 3297 19150 3303 19167
rect 3320 19166 3326 19167
rect 3549 19166 3552 19172
rect 3320 19152 3552 19166
rect 3320 19150 3326 19152
rect 3297 19147 3326 19150
rect 3549 19146 3552 19152
rect 3578 19146 3581 19172
rect 5573 19146 5576 19172
rect 5602 19166 5605 19172
rect 6962 19170 6976 19254
rect 8241 19248 8244 19254
rect 8270 19248 8273 19274
rect 8449 19269 8478 19272
rect 8449 19252 8455 19269
rect 8472 19268 8478 19269
rect 8839 19268 8842 19274
rect 8472 19254 8842 19268
rect 8472 19252 8478 19254
rect 8449 19249 8478 19252
rect 8839 19248 8842 19254
rect 8868 19248 8871 19274
rect 17717 19248 17720 19274
rect 17746 19268 17749 19274
rect 19235 19268 19238 19274
rect 17746 19254 19238 19268
rect 17746 19248 17749 19254
rect 7275 19180 7278 19206
rect 7304 19200 7307 19206
rect 18922 19204 18936 19254
rect 19235 19248 19238 19254
rect 19264 19268 19267 19274
rect 19327 19268 19330 19274
rect 19264 19254 19330 19268
rect 19264 19248 19267 19254
rect 19327 19248 19330 19254
rect 19356 19248 19359 19274
rect 19949 19269 19978 19272
rect 19949 19252 19955 19269
rect 19972 19268 19978 19269
rect 20293 19268 20296 19274
rect 19972 19254 20296 19268
rect 19972 19252 19978 19254
rect 19949 19249 19978 19252
rect 20293 19248 20296 19254
rect 20322 19248 20325 19274
rect 22479 19269 22508 19272
rect 22479 19252 22485 19269
rect 22502 19268 22508 19269
rect 22777 19268 22780 19274
rect 22502 19254 22780 19268
rect 22502 19252 22508 19254
rect 22479 19249 22508 19252
rect 22777 19248 22780 19254
rect 22806 19248 22809 19274
rect 25537 19248 25540 19274
rect 25566 19268 25569 19274
rect 25629 19268 25632 19274
rect 25566 19254 25632 19268
rect 25566 19248 25569 19254
rect 25629 19248 25632 19254
rect 25658 19248 25661 19274
rect 26687 19214 26690 19240
rect 26716 19234 26719 19240
rect 27240 19235 27269 19238
rect 27240 19234 27246 19235
rect 26716 19220 27246 19234
rect 26716 19214 26719 19220
rect 27240 19218 27246 19220
rect 27263 19218 27269 19235
rect 27240 19215 27269 19218
rect 7414 19201 7443 19204
rect 7414 19200 7420 19201
rect 7304 19186 7420 19200
rect 7304 19180 7307 19186
rect 7414 19184 7420 19186
rect 7437 19184 7443 19201
rect 7414 19181 7443 19184
rect 18914 19201 18943 19204
rect 18914 19184 18920 19201
rect 18937 19184 18943 19201
rect 18914 19181 18943 19184
rect 20707 19180 20710 19206
rect 20736 19200 20739 19206
rect 20736 19186 21512 19200
rect 20736 19180 20739 19186
rect 6954 19167 6983 19170
rect 5602 19152 5760 19166
rect 5602 19146 5605 19152
rect 3365 19136 3368 19138
rect 3347 19133 3368 19136
rect 3347 19116 3353 19133
rect 3347 19113 3368 19116
rect 3365 19112 3368 19113
rect 3394 19112 3397 19138
rect 5746 19136 5760 19152
rect 6954 19150 6960 19167
rect 6977 19150 6983 19167
rect 6954 19147 6983 19150
rect 7613 19167 7642 19170
rect 7613 19150 7619 19167
rect 7636 19166 7642 19167
rect 8287 19166 8290 19172
rect 7636 19152 8290 19166
rect 7636 19150 7642 19152
rect 7613 19147 7642 19150
rect 8287 19146 8290 19152
rect 8316 19166 8319 19172
rect 8471 19166 8474 19172
rect 8316 19152 8474 19166
rect 8316 19146 8319 19152
rect 8471 19146 8474 19152
rect 8500 19146 8503 19172
rect 18637 19146 18640 19172
rect 18666 19166 18669 19172
rect 19113 19167 19142 19170
rect 19113 19166 19119 19167
rect 18666 19152 19119 19166
rect 18666 19146 18669 19152
rect 19113 19150 19119 19152
rect 19136 19150 19142 19167
rect 19113 19147 19142 19150
rect 21259 19146 21262 19172
rect 21288 19166 21291 19172
rect 21351 19166 21354 19172
rect 21288 19152 21354 19166
rect 21288 19146 21291 19152
rect 21351 19146 21354 19152
rect 21380 19166 21383 19172
rect 21444 19167 21473 19170
rect 21444 19166 21450 19167
rect 21380 19152 21450 19166
rect 21380 19146 21383 19152
rect 21444 19150 21450 19152
rect 21467 19150 21473 19167
rect 21498 19166 21512 19186
rect 24350 19186 24456 19200
rect 21643 19167 21672 19170
rect 21643 19166 21649 19167
rect 21498 19152 21649 19166
rect 21444 19147 21473 19150
rect 21643 19150 21649 19152
rect 21666 19166 21672 19167
rect 24350 19166 24364 19186
rect 21666 19152 24364 19166
rect 24388 19167 24417 19170
rect 21666 19150 21672 19152
rect 21643 19147 21672 19150
rect 24388 19150 24394 19167
rect 24411 19150 24417 19167
rect 24442 19166 24456 19186
rect 27377 19180 27380 19206
rect 27406 19180 27409 19206
rect 24587 19167 24616 19170
rect 24587 19166 24593 19167
rect 24442 19152 24593 19166
rect 24388 19147 24417 19150
rect 24587 19150 24593 19152
rect 24610 19166 24616 19167
rect 27194 19167 27223 19170
rect 24610 19152 25537 19166
rect 24610 19150 24616 19152
rect 24587 19147 24616 19150
rect 5688 19133 5717 19136
rect 5688 19132 5694 19133
rect 5582 19118 5694 19132
rect 5582 19104 5596 19118
rect 5688 19116 5694 19118
rect 5711 19116 5717 19133
rect 5688 19113 5717 19116
rect 5739 19133 5768 19136
rect 5739 19116 5745 19133
rect 5762 19116 5768 19133
rect 5739 19113 5768 19116
rect 6815 19112 6818 19138
rect 6844 19112 6847 19138
rect 6907 19112 6910 19138
rect 6936 19112 6939 19138
rect 7413 19112 7416 19138
rect 7442 19132 7445 19138
rect 7574 19133 7603 19136
rect 7574 19132 7580 19133
rect 7442 19118 7580 19132
rect 7442 19112 7445 19118
rect 7574 19116 7580 19118
rect 7597 19116 7603 19133
rect 19074 19133 19103 19136
rect 19074 19132 19080 19133
rect 7574 19113 7603 19116
rect 18968 19118 19080 19132
rect 5573 19078 5576 19104
rect 5602 19078 5605 19104
rect 6539 19078 6542 19104
rect 6568 19102 6571 19104
rect 6568 19099 6592 19102
rect 6568 19082 6569 19099
rect 6586 19082 6592 19099
rect 6568 19079 6592 19082
rect 6568 19078 6571 19079
rect 12105 19078 12108 19104
rect 12134 19098 12137 19104
rect 12979 19098 12982 19104
rect 12134 19084 12982 19098
rect 12134 19078 12137 19084
rect 12979 19078 12982 19084
rect 13008 19078 13011 19104
rect 17947 19078 17950 19104
rect 17976 19098 17979 19104
rect 18968 19098 18982 19118
rect 19074 19116 19080 19118
rect 19097 19116 19103 19133
rect 19074 19113 19103 19116
rect 21029 19112 21032 19138
rect 21058 19132 21061 19138
rect 21604 19133 21633 19136
rect 21604 19132 21610 19133
rect 21058 19118 21610 19132
rect 21058 19112 21061 19118
rect 21604 19116 21610 19118
rect 21627 19116 21633 19133
rect 21604 19113 21633 19116
rect 17976 19084 18982 19098
rect 17976 19078 17979 19084
rect 24157 19078 24160 19104
rect 24186 19098 24189 19104
rect 24396 19098 24410 19147
rect 24433 19112 24436 19138
rect 24462 19132 24465 19138
rect 24548 19133 24577 19136
rect 24548 19132 24554 19133
rect 24462 19118 24554 19132
rect 24462 19112 24465 19118
rect 24548 19116 24554 19118
rect 24571 19116 24577 19133
rect 25523 19132 25537 19152
rect 27194 19150 27200 19167
rect 27217 19166 27223 19167
rect 29539 19166 29542 19172
rect 27217 19152 29542 19166
rect 27217 19150 27223 19152
rect 27194 19147 27223 19150
rect 29539 19146 29542 19152
rect 29568 19146 29571 19172
rect 28619 19132 28622 19138
rect 25523 19118 28622 19132
rect 24548 19113 24577 19116
rect 28619 19112 28622 19118
rect 28648 19112 28651 19138
rect 24186 19084 24410 19098
rect 25423 19099 25452 19102
rect 24186 19078 24189 19084
rect 25423 19082 25429 19099
rect 25446 19098 25452 19099
rect 25491 19098 25494 19104
rect 25446 19084 25494 19098
rect 25446 19082 25452 19084
rect 25423 19079 25452 19082
rect 25491 19078 25494 19084
rect 25520 19078 25523 19104
rect 27239 19078 27242 19104
rect 27268 19078 27271 19104
rect 27285 19078 27288 19104
rect 27314 19078 27317 19104
rect 3036 19016 29992 19064
rect 4837 18976 4840 19002
rect 4866 18976 4869 19002
rect 6448 18997 6477 19000
rect 6448 18980 6454 18997
rect 6471 18996 6477 18997
rect 6815 18996 6818 19002
rect 6471 18982 6818 18996
rect 6471 18980 6477 18982
rect 6448 18977 6477 18980
rect 6815 18976 6818 18982
rect 6844 18976 6847 19002
rect 8311 18997 8340 19000
rect 8311 18980 8317 18997
rect 8334 18996 8340 18997
rect 8977 18996 8980 19002
rect 8334 18982 8980 18996
rect 8334 18980 8340 18982
rect 8311 18977 8340 18980
rect 8977 18976 8980 18982
rect 9006 18976 9009 19002
rect 14957 18976 14960 19002
rect 14986 18996 14989 19002
rect 14986 18982 15348 18996
rect 14986 18976 14989 18982
rect 3623 18963 3652 18966
rect 3623 18946 3629 18963
rect 3646 18962 3652 18963
rect 3687 18962 3690 18968
rect 3646 18948 3690 18962
rect 3646 18946 3652 18948
rect 3623 18943 3652 18946
rect 3687 18942 3690 18948
rect 3716 18942 3719 18968
rect 4700 18963 4729 18966
rect 4700 18946 4706 18963
rect 4723 18962 4729 18963
rect 4846 18962 4860 18976
rect 4723 18948 4860 18962
rect 4723 18946 4729 18948
rect 4700 18943 4729 18946
rect 6493 18942 6496 18968
rect 6522 18942 6525 18968
rect 6539 18942 6542 18968
rect 6568 18942 6571 18968
rect 7505 18966 7508 18968
rect 7487 18963 7508 18966
rect 7487 18946 7493 18963
rect 7487 18943 7508 18946
rect 7505 18942 7508 18943
rect 7534 18942 7537 18968
rect 12041 18963 12070 18966
rect 12041 18946 12047 18963
rect 12064 18962 12070 18963
rect 12064 18948 12174 18962
rect 12064 18946 12070 18948
rect 12041 18943 12070 18946
rect 3135 18908 3138 18934
rect 3164 18928 3167 18934
rect 3412 18929 3441 18932
rect 3412 18928 3418 18929
rect 3164 18914 3418 18928
rect 3164 18908 3167 18914
rect 3412 18912 3418 18914
rect 3435 18912 3441 18929
rect 3412 18909 3441 18912
rect 3549 18908 3552 18934
rect 3578 18932 3581 18934
rect 3578 18929 3596 18932
rect 3590 18912 3596 18929
rect 3578 18909 3596 18912
rect 4792 18929 4821 18932
rect 4792 18912 4798 18929
rect 4815 18912 4821 18929
rect 4792 18909 4821 18912
rect 3578 18908 3581 18909
rect 4699 18874 4702 18900
rect 4728 18894 4731 18900
rect 4800 18894 4814 18909
rect 4837 18908 4840 18934
rect 4866 18908 4869 18934
rect 6356 18929 6385 18932
rect 6356 18928 6362 18929
rect 6203 18914 6362 18928
rect 4728 18880 4814 18894
rect 4728 18874 4731 18880
rect 4838 18861 4867 18864
rect 4838 18844 4844 18861
rect 4861 18860 4867 18861
rect 6203 18860 6217 18914
rect 6356 18912 6362 18914
rect 6379 18912 6385 18929
rect 6356 18909 6385 18912
rect 6401 18908 6404 18934
rect 6430 18908 6433 18934
rect 6586 18929 6615 18932
rect 6586 18912 6592 18929
rect 6609 18928 6615 18929
rect 6631 18928 6634 18934
rect 6609 18914 6634 18928
rect 6609 18912 6615 18914
rect 6586 18909 6615 18912
rect 6631 18908 6634 18914
rect 6660 18908 6663 18934
rect 7275 18908 7278 18934
rect 7304 18908 7307 18934
rect 7413 18928 7416 18934
rect 7442 18932 7445 18934
rect 7442 18929 7460 18932
rect 7330 18914 7416 18928
rect 6953 18874 6956 18900
rect 6982 18894 6985 18900
rect 7330 18894 7344 18914
rect 7413 18908 7416 18914
rect 7454 18912 7460 18929
rect 7442 18909 7460 18912
rect 7442 18908 7445 18909
rect 11461 18908 11464 18934
rect 11490 18928 11493 18934
rect 11985 18929 12014 18932
rect 11985 18928 11991 18929
rect 11490 18914 11991 18928
rect 11490 18908 11493 18914
rect 11985 18912 11991 18914
rect 12008 18928 12014 18929
rect 12105 18928 12108 18934
rect 12008 18914 12108 18928
rect 12008 18912 12014 18914
rect 11985 18909 12014 18912
rect 12105 18908 12108 18914
rect 12134 18908 12137 18934
rect 12160 18928 12174 18948
rect 14313 18942 14316 18968
rect 14342 18962 14345 18968
rect 14474 18963 14503 18966
rect 14474 18962 14480 18963
rect 14342 18948 14480 18962
rect 14342 18942 14345 18948
rect 14474 18946 14480 18948
rect 14497 18946 14503 18963
rect 14474 18943 14503 18946
rect 14525 18963 14554 18966
rect 14525 18946 14531 18963
rect 14548 18962 14554 18963
rect 15334 18962 15348 18982
rect 24295 18976 24298 19002
rect 24324 18996 24327 19002
rect 24388 18997 24417 19000
rect 24388 18996 24394 18997
rect 24324 18982 24394 18996
rect 24324 18976 24327 18982
rect 24388 18980 24394 18982
rect 24411 18980 24417 18997
rect 24388 18977 24417 18980
rect 24663 18976 24666 19002
rect 24692 18996 24695 19002
rect 24756 18997 24785 19000
rect 24756 18996 24762 18997
rect 24692 18982 24762 18996
rect 24692 18976 24695 18982
rect 24756 18980 24762 18982
rect 24779 18980 24785 18997
rect 24756 18977 24785 18980
rect 24802 18997 24831 19000
rect 24802 18980 24808 18997
rect 24825 18996 24831 18997
rect 24825 18982 25422 18996
rect 24825 18980 24831 18982
rect 24802 18977 24831 18980
rect 17883 18963 17912 18966
rect 14548 18946 14566 18962
rect 15334 18948 15670 18962
rect 14525 18943 14566 18946
rect 12427 18928 12430 18934
rect 12160 18914 12430 18928
rect 12427 18908 12430 18914
rect 12456 18928 12459 18934
rect 12565 18928 12568 18934
rect 12456 18914 12568 18928
rect 12456 18908 12459 18914
rect 12565 18908 12568 18914
rect 12594 18908 12597 18934
rect 14552 18928 14566 18943
rect 14589 18928 14592 18934
rect 14552 18914 14592 18928
rect 14589 18908 14592 18914
rect 14618 18928 14621 18934
rect 15049 18928 15052 18934
rect 14618 18914 15052 18928
rect 14618 18908 14621 18914
rect 15049 18908 15052 18914
rect 15078 18908 15081 18934
rect 15349 18929 15378 18932
rect 15349 18912 15355 18929
rect 15372 18928 15378 18929
rect 15602 18929 15631 18932
rect 15602 18928 15608 18929
rect 15372 18914 15608 18928
rect 15372 18912 15378 18914
rect 15349 18909 15378 18912
rect 15602 18912 15608 18914
rect 15625 18912 15631 18929
rect 15656 18928 15670 18948
rect 17883 18946 17889 18963
rect 17906 18962 17912 18963
rect 17906 18948 18016 18962
rect 17906 18946 17912 18948
rect 17883 18943 17912 18946
rect 15693 18928 15696 18934
rect 15656 18914 15696 18928
rect 15602 18909 15631 18912
rect 15693 18908 15696 18914
rect 15722 18908 15725 18934
rect 15739 18908 15742 18934
rect 15768 18908 15771 18934
rect 15789 18929 15818 18932
rect 15789 18912 15795 18929
rect 15812 18912 15818 18929
rect 15789 18909 15818 18912
rect 17672 18929 17701 18932
rect 17672 18912 17678 18929
rect 17695 18928 17701 18929
rect 17717 18928 17720 18934
rect 17695 18914 17720 18928
rect 17695 18912 17701 18914
rect 17672 18909 17701 18912
rect 6982 18880 7344 18894
rect 6982 18874 6985 18880
rect 11829 18874 11832 18900
rect 11858 18874 11861 18900
rect 14083 18874 14086 18900
rect 14112 18894 14115 18900
rect 14314 18895 14343 18898
rect 14314 18894 14320 18895
rect 14112 18880 14320 18894
rect 14112 18874 14115 18880
rect 14314 18878 14320 18880
rect 14337 18878 14343 18895
rect 14314 18875 14343 18878
rect 15279 18874 15282 18900
rect 15308 18894 15311 18900
rect 15647 18894 15650 18900
rect 15308 18880 15650 18894
rect 15308 18874 15311 18880
rect 15647 18874 15650 18880
rect 15676 18894 15679 18900
rect 15794 18894 15808 18909
rect 17717 18908 17720 18914
rect 17746 18908 17749 18934
rect 17833 18929 17862 18932
rect 17833 18912 17839 18929
rect 17856 18928 17862 18929
rect 17947 18928 17950 18934
rect 17856 18914 17950 18928
rect 17856 18912 17862 18914
rect 17833 18909 17862 18912
rect 17947 18908 17950 18914
rect 17976 18908 17979 18934
rect 18002 18928 18016 18948
rect 21351 18942 21354 18968
rect 21380 18962 21383 18968
rect 22961 18962 22964 18968
rect 21380 18948 22964 18962
rect 21380 18942 21383 18948
rect 22961 18942 22964 18948
rect 22990 18942 22993 18968
rect 23127 18963 23156 18966
rect 23127 18946 23133 18963
rect 23150 18962 23156 18963
rect 23150 18948 23260 18962
rect 23150 18946 23156 18948
rect 23127 18943 23156 18946
rect 20707 18928 20710 18934
rect 18002 18914 20710 18928
rect 20707 18908 20710 18914
rect 20736 18908 20739 18934
rect 15676 18880 15808 18894
rect 22916 18895 22945 18898
rect 15676 18874 15679 18880
rect 22916 18878 22922 18895
rect 22939 18894 22945 18895
rect 22970 18894 22984 18942
rect 23246 18934 23260 18948
rect 24111 18942 24114 18968
rect 24140 18962 24143 18968
rect 24433 18962 24436 18968
rect 24140 18948 24436 18962
rect 24140 18942 24143 18948
rect 24433 18942 24436 18948
rect 24462 18942 24465 18968
rect 23077 18929 23106 18932
rect 23077 18912 23083 18929
rect 23100 18928 23106 18929
rect 23191 18928 23194 18934
rect 23100 18914 23194 18928
rect 23100 18912 23106 18914
rect 23077 18909 23106 18912
rect 23191 18908 23194 18914
rect 23220 18908 23223 18934
rect 23237 18908 23240 18934
rect 23266 18908 23269 18934
rect 24249 18908 24252 18934
rect 24278 18928 24281 18934
rect 24296 18929 24325 18932
rect 24296 18928 24302 18929
rect 24278 18914 24302 18928
rect 24278 18908 24281 18914
rect 24296 18912 24302 18914
rect 24319 18912 24325 18929
rect 24296 18909 24325 18912
rect 24341 18908 24344 18934
rect 24370 18908 24373 18934
rect 24480 18929 24509 18932
rect 24480 18912 24486 18929
rect 24503 18928 24509 18929
rect 24710 18929 24739 18932
rect 24710 18928 24716 18929
rect 24503 18914 24716 18928
rect 24503 18912 24509 18914
rect 24480 18909 24509 18912
rect 24710 18912 24716 18914
rect 24733 18912 24739 18929
rect 24710 18909 24739 18912
rect 25353 18908 25356 18934
rect 25382 18908 25385 18934
rect 25408 18898 25422 18982
rect 25491 18942 25494 18968
rect 25520 18942 25523 18968
rect 26503 18966 26506 18968
rect 26485 18963 26506 18966
rect 26485 18946 26491 18963
rect 26485 18943 26506 18946
rect 26503 18942 26506 18943
rect 26532 18942 26535 18968
rect 28417 18963 28446 18966
rect 28417 18946 28423 18963
rect 28440 18962 28446 18963
rect 28440 18948 28550 18962
rect 28440 18946 28446 18948
rect 28417 18943 28446 18946
rect 28536 18934 28550 18948
rect 25445 18908 25448 18934
rect 25474 18908 25477 18934
rect 25541 18924 25570 18927
rect 25541 18907 25547 18924
rect 25564 18907 25570 18924
rect 25629 18908 25632 18934
rect 25658 18928 25661 18934
rect 25721 18928 25724 18934
rect 25658 18914 25724 18928
rect 25658 18908 25661 18914
rect 25721 18908 25724 18914
rect 25750 18928 25753 18934
rect 26429 18929 26458 18932
rect 26429 18928 26435 18929
rect 25750 18914 26435 18928
rect 25750 18908 25753 18914
rect 26429 18912 26435 18914
rect 26452 18912 26458 18929
rect 26429 18909 26458 18912
rect 28021 18908 28024 18934
rect 28050 18928 28053 18934
rect 28206 18929 28235 18932
rect 28206 18928 28212 18929
rect 28050 18914 28212 18928
rect 28050 18908 28053 18914
rect 28206 18912 28212 18914
rect 28229 18912 28235 18929
rect 28206 18909 28235 18912
rect 28343 18908 28346 18934
rect 28372 18932 28375 18934
rect 28372 18929 28390 18932
rect 28384 18912 28390 18929
rect 28372 18909 28390 18912
rect 28372 18908 28375 18909
rect 28527 18908 28530 18934
rect 28556 18908 28559 18934
rect 29241 18929 29270 18932
rect 29241 18912 29247 18929
rect 29264 18928 29270 18929
rect 29494 18929 29523 18932
rect 29494 18928 29500 18929
rect 29264 18914 29500 18928
rect 29264 18912 29270 18914
rect 29241 18909 29270 18912
rect 29494 18912 29500 18914
rect 29517 18912 29523 18929
rect 29494 18909 29523 18912
rect 29585 18908 29588 18934
rect 29614 18908 29617 18934
rect 29631 18908 29634 18934
rect 29660 18908 29663 18934
rect 29677 18908 29680 18934
rect 29706 18932 29709 18934
rect 29706 18909 29710 18932
rect 29706 18908 29709 18909
rect 25541 18904 25570 18907
rect 24894 18895 24923 18898
rect 22939 18880 22984 18894
rect 23890 18880 24824 18894
rect 22939 18878 22945 18880
rect 22916 18875 22945 18878
rect 4861 18846 6217 18860
rect 4861 18844 4867 18846
rect 4838 18841 4867 18844
rect 4447 18827 4476 18830
rect 4447 18810 4453 18827
rect 4470 18826 4476 18827
rect 4975 18826 4978 18832
rect 4470 18812 4978 18826
rect 4470 18810 4476 18812
rect 4447 18807 4476 18810
rect 4975 18806 4978 18812
rect 5004 18806 5007 18832
rect 8563 18806 8566 18832
rect 8592 18826 8595 18832
rect 9069 18826 9072 18832
rect 8592 18812 9072 18826
rect 8592 18806 8595 18812
rect 9069 18806 9072 18812
rect 9098 18826 9101 18832
rect 9529 18826 9532 18832
rect 9098 18812 9532 18826
rect 9098 18806 9101 18812
rect 9529 18806 9532 18812
rect 9558 18806 9561 18832
rect 12865 18827 12894 18830
rect 12865 18810 12871 18827
rect 12888 18826 12894 18827
rect 13071 18826 13074 18832
rect 12888 18812 13074 18826
rect 12888 18810 12894 18812
rect 12865 18807 12894 18810
rect 13071 18806 13074 18812
rect 13100 18806 13103 18832
rect 15602 18827 15631 18830
rect 15602 18810 15608 18827
rect 15625 18826 15631 18827
rect 15693 18826 15696 18832
rect 15625 18812 15696 18826
rect 15625 18810 15631 18812
rect 15602 18807 15631 18810
rect 15693 18806 15696 18812
rect 15722 18806 15725 18832
rect 18707 18827 18736 18830
rect 18707 18810 18713 18827
rect 18730 18826 18736 18827
rect 19143 18826 19146 18832
rect 18730 18812 19146 18826
rect 18730 18810 18736 18812
rect 18707 18807 18736 18810
rect 19143 18806 19146 18812
rect 19172 18806 19175 18832
rect 22915 18806 22918 18832
rect 22944 18826 22947 18832
rect 23890 18826 23904 18880
rect 24019 18840 24022 18866
rect 24048 18860 24051 18866
rect 24204 18861 24233 18864
rect 24204 18860 24210 18861
rect 24048 18846 24210 18860
rect 24048 18840 24051 18846
rect 24204 18844 24210 18846
rect 24227 18844 24233 18861
rect 24204 18841 24233 18844
rect 22944 18812 23904 18826
rect 23951 18827 23980 18830
rect 22944 18806 22947 18812
rect 23951 18810 23957 18827
rect 23974 18826 23980 18827
rect 24295 18826 24298 18832
rect 23974 18812 24298 18826
rect 23974 18810 23980 18812
rect 23951 18807 23980 18810
rect 24295 18806 24298 18812
rect 24324 18806 24327 18832
rect 24663 18806 24666 18832
rect 24692 18826 24695 18832
rect 24756 18827 24785 18830
rect 24756 18826 24762 18827
rect 24692 18812 24762 18826
rect 24692 18806 24695 18812
rect 24756 18810 24762 18812
rect 24779 18810 24785 18827
rect 24810 18826 24824 18880
rect 24894 18878 24900 18895
rect 24917 18878 24923 18895
rect 24894 18875 24923 18878
rect 25400 18895 25429 18898
rect 25400 18878 25406 18895
rect 25423 18878 25429 18895
rect 25400 18875 25429 18878
rect 24902 18860 24916 18875
rect 25491 18860 25494 18866
rect 24902 18846 25494 18860
rect 25491 18840 25494 18846
rect 25520 18840 25523 18866
rect 25546 18826 25560 18904
rect 26274 18895 26303 18898
rect 26274 18878 26280 18895
rect 26297 18878 26303 18895
rect 26274 18875 26303 18878
rect 24810 18812 25560 18826
rect 26282 18826 26296 18875
rect 29539 18874 29542 18900
rect 29568 18874 29571 18900
rect 27975 18860 27978 18866
rect 27110 18846 27978 18860
rect 27110 18826 27124 18846
rect 27975 18840 27978 18846
rect 28004 18840 28007 18866
rect 26282 18812 27124 18826
rect 27309 18827 27338 18830
rect 24756 18807 24785 18810
rect 27309 18810 27315 18827
rect 27332 18826 27338 18827
rect 27377 18826 27380 18832
rect 27332 18812 27380 18826
rect 27332 18810 27338 18812
rect 27309 18807 27338 18810
rect 27377 18806 27380 18812
rect 27406 18806 27409 18832
rect 3036 18744 29992 18792
rect 4654 18725 4683 18728
rect 4654 18708 4660 18725
rect 4677 18724 4683 18725
rect 4837 18724 4840 18730
rect 4677 18710 4840 18724
rect 4677 18708 4683 18710
rect 4654 18705 4683 18708
rect 4837 18704 4840 18710
rect 4866 18704 4869 18730
rect 5665 18724 5668 18730
rect 5260 18710 5668 18724
rect 4856 18623 4885 18626
rect 4856 18606 4862 18623
rect 4879 18622 4885 18623
rect 5067 18622 5070 18628
rect 4879 18608 5070 18622
rect 4879 18606 4885 18608
rect 4856 18603 4885 18606
rect 5067 18602 5070 18608
rect 5096 18602 5099 18628
rect 5260 18626 5274 18710
rect 5665 18704 5668 18710
rect 5694 18704 5697 18730
rect 10357 18704 10360 18730
rect 10386 18724 10389 18730
rect 10864 18725 10893 18728
rect 10864 18724 10870 18725
rect 10386 18710 10870 18724
rect 10386 18704 10389 18710
rect 10864 18708 10870 18710
rect 10887 18708 10893 18725
rect 10864 18705 10893 18708
rect 15211 18725 15240 18728
rect 15211 18708 15217 18725
rect 15234 18724 15240 18725
rect 15739 18724 15742 18730
rect 15234 18710 15742 18724
rect 15234 18708 15240 18710
rect 15211 18705 15240 18708
rect 15739 18704 15742 18710
rect 15768 18704 15771 18730
rect 22593 18724 22596 18730
rect 22096 18710 22596 18724
rect 12979 18670 12982 18696
rect 13008 18690 13011 18696
rect 20524 18691 20553 18694
rect 13008 18676 14198 18690
rect 13008 18670 13011 18676
rect 13026 18657 13055 18660
rect 13026 18640 13032 18657
rect 13049 18656 13055 18657
rect 13669 18656 13672 18662
rect 13049 18642 13672 18656
rect 13049 18640 13055 18642
rect 13026 18637 13055 18640
rect 13669 18636 13672 18642
rect 13698 18636 13701 18662
rect 14184 18656 14198 18676
rect 15610 18676 15877 18690
rect 15141 18656 15144 18662
rect 14184 18642 14244 18656
rect 5252 18623 5281 18626
rect 5252 18606 5258 18623
rect 5275 18606 5281 18623
rect 5252 18603 5281 18606
rect 5413 18623 5442 18626
rect 5413 18606 5419 18623
rect 5436 18622 5442 18623
rect 5803 18622 5806 18628
rect 5436 18608 5806 18622
rect 5436 18606 5442 18608
rect 5413 18603 5442 18606
rect 5803 18602 5806 18608
rect 5832 18602 5835 18628
rect 8287 18602 8290 18628
rect 8316 18602 8319 18628
rect 8449 18623 8478 18626
rect 8449 18606 8455 18623
rect 8472 18622 8478 18623
rect 8563 18622 8566 18628
rect 8472 18608 8566 18622
rect 8472 18606 8478 18608
rect 8449 18603 8478 18606
rect 8563 18602 8566 18608
rect 8592 18602 8595 18628
rect 9345 18622 9348 18628
rect 8618 18608 9348 18622
rect 4653 18568 4656 18594
rect 4682 18568 4685 18594
rect 4746 18589 4775 18592
rect 4746 18572 4752 18589
rect 4769 18572 4775 18589
rect 4746 18569 4775 18572
rect 4754 18554 4768 18569
rect 4791 18568 4794 18594
rect 4820 18568 4823 18594
rect 5481 18592 5484 18594
rect 5463 18589 5484 18592
rect 5463 18588 5469 18589
rect 5260 18574 5469 18588
rect 5260 18560 5274 18574
rect 5463 18572 5469 18574
rect 5463 18569 5484 18572
rect 5481 18568 5484 18569
rect 5510 18568 5513 18594
rect 8517 18592 8520 18594
rect 8499 18589 8520 18592
rect 8499 18572 8505 18589
rect 8546 18588 8549 18594
rect 8618 18588 8632 18608
rect 9345 18602 9348 18608
rect 9374 18602 9377 18628
rect 10771 18602 10774 18628
rect 10800 18622 10803 18628
rect 10956 18623 10985 18626
rect 10956 18622 10962 18623
rect 10800 18608 10962 18622
rect 10800 18602 10803 18608
rect 10956 18606 10962 18608
rect 10979 18606 10985 18623
rect 10956 18603 10985 18606
rect 11047 18602 11050 18628
rect 11076 18626 11079 18628
rect 11076 18603 11080 18626
rect 11416 18623 11445 18626
rect 11416 18606 11422 18623
rect 11439 18622 11445 18623
rect 11829 18622 11832 18628
rect 11439 18608 11832 18622
rect 11439 18606 11445 18608
rect 11416 18603 11445 18606
rect 11076 18602 11079 18603
rect 8546 18574 8632 18588
rect 8499 18569 8520 18572
rect 8517 18568 8520 18569
rect 8546 18568 8549 18574
rect 10863 18568 10866 18594
rect 10892 18568 10895 18594
rect 11001 18568 11004 18594
rect 11030 18568 11033 18594
rect 5113 18554 5116 18560
rect 4754 18540 5116 18554
rect 5113 18534 5116 18540
rect 5142 18534 5145 18560
rect 5251 18534 5254 18560
rect 5280 18534 5283 18560
rect 6263 18534 6266 18560
rect 6292 18558 6295 18560
rect 6292 18555 6316 18558
rect 6292 18538 6293 18555
rect 6310 18538 6316 18555
rect 6292 18535 6316 18538
rect 9323 18555 9352 18558
rect 9323 18538 9329 18555
rect 9346 18554 9352 18555
rect 9483 18554 9486 18560
rect 9346 18540 9486 18554
rect 9346 18538 9352 18540
rect 9323 18535 9352 18538
rect 6292 18534 6295 18535
rect 9483 18534 9486 18540
rect 9512 18534 9515 18560
rect 10909 18534 10912 18560
rect 10938 18554 10941 18560
rect 11424 18554 11438 18603
rect 11829 18602 11832 18608
rect 11858 18602 11861 18628
rect 13071 18602 13074 18628
rect 13100 18602 13103 18628
rect 13117 18602 13120 18628
rect 13146 18626 13149 18628
rect 13146 18622 13150 18626
rect 13146 18608 13168 18622
rect 13146 18603 13150 18608
rect 13146 18602 13149 18603
rect 13853 18602 13856 18628
rect 13882 18622 13885 18628
rect 14083 18622 14086 18628
rect 13882 18608 14086 18622
rect 13882 18602 13885 18608
rect 14083 18602 14086 18608
rect 14112 18622 14115 18628
rect 14176 18623 14205 18626
rect 14176 18622 14182 18623
rect 14112 18608 14182 18622
rect 14112 18602 14115 18608
rect 14176 18606 14182 18608
rect 14199 18606 14205 18623
rect 14230 18622 14244 18642
rect 15058 18642 15144 18656
rect 15058 18628 15072 18642
rect 15141 18636 15144 18642
rect 15170 18636 15173 18662
rect 14313 18622 14316 18628
rect 14342 18626 14345 18628
rect 14342 18623 14360 18626
rect 14230 18608 14316 18622
rect 14176 18603 14205 18606
rect 14313 18602 14316 18608
rect 14354 18622 14360 18623
rect 15049 18622 15052 18628
rect 14354 18608 15052 18622
rect 14354 18606 14360 18608
rect 14342 18603 14360 18606
rect 14342 18602 14345 18603
rect 15049 18602 15052 18608
rect 15078 18622 15081 18628
rect 15610 18622 15624 18676
rect 15647 18636 15650 18662
rect 15676 18656 15679 18662
rect 15785 18656 15788 18662
rect 15676 18642 15788 18656
rect 15676 18636 15679 18642
rect 15785 18636 15788 18642
rect 15814 18636 15817 18662
rect 15863 18656 15877 18676
rect 20524 18674 20530 18691
rect 20547 18690 20553 18691
rect 20547 18676 21328 18690
rect 20547 18674 20553 18676
rect 20524 18671 20553 18674
rect 15863 18642 15946 18656
rect 15078 18608 15624 18622
rect 15078 18602 15081 18608
rect 15693 18602 15696 18628
rect 15722 18602 15725 18628
rect 15878 18623 15907 18626
rect 15878 18606 15884 18623
rect 15901 18606 15907 18623
rect 15878 18603 15907 18606
rect 11461 18568 11464 18594
rect 11490 18588 11493 18594
rect 11645 18592 11648 18594
rect 11576 18589 11605 18592
rect 11576 18588 11582 18589
rect 11490 18574 11582 18588
rect 11490 18568 11493 18574
rect 11576 18572 11582 18574
rect 11599 18572 11605 18589
rect 11576 18569 11605 18572
rect 11627 18589 11648 18592
rect 11627 18572 11633 18589
rect 11627 18569 11648 18572
rect 11645 18568 11648 18569
rect 11674 18568 11677 18594
rect 12451 18589 12480 18592
rect 12451 18572 12457 18589
rect 12474 18588 12480 18589
rect 12934 18589 12963 18592
rect 12934 18588 12940 18589
rect 12474 18574 12940 18588
rect 12474 18572 12480 18574
rect 12451 18569 12480 18572
rect 12934 18572 12940 18574
rect 12957 18572 12963 18589
rect 12934 18569 12963 18572
rect 13026 18589 13055 18592
rect 13026 18572 13032 18589
rect 13049 18572 13055 18589
rect 13026 18569 13055 18572
rect 14387 18589 14416 18592
rect 14387 18572 14393 18589
rect 14410 18588 14416 18589
rect 14451 18588 14454 18594
rect 14410 18574 14454 18588
rect 14410 18572 14416 18574
rect 14387 18569 14416 18572
rect 10938 18540 11438 18554
rect 13034 18554 13048 18569
rect 14451 18568 14454 18574
rect 14480 18568 14483 18594
rect 15233 18568 15236 18594
rect 15262 18588 15265 18594
rect 15886 18588 15900 18603
rect 15262 18574 15900 18588
rect 15932 18588 15946 18642
rect 18453 18636 18456 18662
rect 18482 18656 18485 18662
rect 18482 18642 19304 18656
rect 18482 18636 18485 18642
rect 15969 18602 15972 18628
rect 15998 18622 16001 18628
rect 16153 18622 16156 18628
rect 15998 18608 16156 18622
rect 15998 18602 16001 18608
rect 16153 18602 16156 18608
rect 16182 18602 16185 18628
rect 16199 18602 16202 18628
rect 16228 18622 16231 18628
rect 16353 18623 16382 18626
rect 16353 18622 16359 18623
rect 16228 18608 16359 18622
rect 16228 18602 16231 18608
rect 16353 18606 16359 18608
rect 16376 18606 16382 18623
rect 16353 18603 16382 18606
rect 19235 18602 19238 18628
rect 19264 18602 19267 18628
rect 19290 18622 19304 18642
rect 20661 18636 20664 18662
rect 20690 18656 20693 18662
rect 20690 18642 20776 18656
rect 20690 18636 20693 18642
rect 19373 18622 19376 18628
rect 19402 18626 19405 18628
rect 19402 18623 19420 18626
rect 19290 18608 19376 18622
rect 19373 18602 19376 18608
rect 19414 18606 19420 18623
rect 20477 18622 20480 18628
rect 19402 18603 19420 18606
rect 19566 18608 20480 18622
rect 19402 18602 19405 18603
rect 16314 18589 16343 18592
rect 16314 18588 16320 18589
rect 15932 18574 16320 18588
rect 15262 18568 15265 18574
rect 16314 18572 16320 18574
rect 16337 18572 16343 18589
rect 16314 18569 16343 18572
rect 19447 18589 19476 18592
rect 19447 18572 19453 18589
rect 19470 18588 19476 18589
rect 19566 18588 19580 18608
rect 20477 18602 20480 18608
rect 20506 18602 20509 18628
rect 20711 18623 20740 18626
rect 20711 18606 20717 18623
rect 20734 18606 20740 18623
rect 20762 18622 20776 18642
rect 21214 18623 21243 18626
rect 21214 18622 21220 18623
rect 20762 18608 21220 18622
rect 20711 18603 20740 18606
rect 21214 18606 21220 18608
rect 21237 18606 21243 18623
rect 21214 18603 21243 18606
rect 19470 18574 19580 18588
rect 20271 18589 20300 18592
rect 19470 18572 19476 18574
rect 19447 18569 19476 18572
rect 20271 18572 20277 18589
rect 20294 18588 20300 18589
rect 20524 18589 20553 18592
rect 20524 18588 20530 18589
rect 20294 18574 20530 18588
rect 20294 18572 20300 18574
rect 20271 18569 20300 18572
rect 20524 18572 20530 18574
rect 20547 18572 20553 18589
rect 20524 18569 20553 18572
rect 20615 18568 20618 18594
rect 20644 18568 20647 18594
rect 20661 18568 20664 18594
rect 20690 18568 20693 18594
rect 20716 18588 20730 18603
rect 20937 18588 20940 18594
rect 20716 18574 20940 18588
rect 20937 18568 20940 18574
rect 20966 18568 20969 18594
rect 13991 18554 13994 18560
rect 13034 18540 13994 18554
rect 10938 18534 10941 18540
rect 13991 18534 13994 18540
rect 14020 18534 14023 18560
rect 15739 18534 15742 18560
rect 15768 18534 15771 18560
rect 15785 18534 15788 18560
rect 15814 18534 15817 18560
rect 15831 18534 15834 18560
rect 15860 18534 15863 18560
rect 17165 18534 17168 18560
rect 17194 18558 17197 18560
rect 17194 18555 17218 18558
rect 17194 18538 17195 18555
rect 17212 18538 17218 18555
rect 17194 18535 17218 18538
rect 17194 18534 17197 18535
rect 21259 18534 21262 18560
rect 21288 18534 21291 18560
rect 21314 18558 21328 18676
rect 22096 18656 22110 18710
rect 22593 18704 22596 18710
rect 22622 18724 22625 18730
rect 25285 18725 25314 18728
rect 22622 18710 25238 18724
rect 22622 18704 22625 18710
rect 22823 18690 22826 18696
rect 22035 18642 22110 18656
rect 22171 18676 22826 18690
rect 21398 18623 21427 18626
rect 21398 18606 21404 18623
rect 21421 18606 21427 18623
rect 21398 18603 21427 18606
rect 21406 18588 21420 18603
rect 21949 18602 21952 18628
rect 21978 18602 21981 18628
rect 22035 18626 22049 18642
rect 22027 18623 22056 18626
rect 22027 18606 22033 18623
rect 22050 18606 22056 18623
rect 22027 18603 22056 18606
rect 22087 18602 22090 18628
rect 22116 18626 22119 18628
rect 22171 18626 22185 18676
rect 22823 18670 22826 18676
rect 22852 18670 22855 18696
rect 25224 18690 25238 18710
rect 25285 18708 25291 18725
rect 25308 18724 25314 18725
rect 25353 18724 25356 18730
rect 25308 18710 25356 18724
rect 25308 18708 25314 18710
rect 25285 18705 25314 18708
rect 25353 18704 25356 18710
rect 25382 18704 25385 18730
rect 27285 18704 27288 18730
rect 27314 18724 27317 18730
rect 27378 18725 27407 18728
rect 27378 18724 27384 18725
rect 27314 18710 27384 18724
rect 27314 18704 27317 18710
rect 27378 18708 27384 18710
rect 27401 18708 27407 18725
rect 27378 18705 27407 18708
rect 25445 18690 25448 18696
rect 25224 18676 25448 18690
rect 25445 18670 25448 18676
rect 25474 18690 25477 18696
rect 27055 18690 27058 18696
rect 25474 18676 27058 18690
rect 25474 18670 25477 18676
rect 27055 18670 27058 18676
rect 27084 18690 27087 18696
rect 27084 18676 27492 18690
rect 27084 18670 27087 18676
rect 22363 18656 22366 18662
rect 22234 18642 22366 18656
rect 22116 18623 22137 18626
rect 22131 18606 22137 18623
rect 22116 18603 22137 18606
rect 22163 18623 22192 18626
rect 22234 18624 22248 18642
rect 22363 18636 22366 18642
rect 22392 18636 22395 18662
rect 24111 18636 24114 18662
rect 24140 18636 24143 18662
rect 26182 18657 26211 18660
rect 26182 18640 26188 18657
rect 26205 18656 26211 18657
rect 26227 18656 26230 18662
rect 26205 18642 26230 18656
rect 26205 18640 26211 18642
rect 26182 18637 26211 18640
rect 26227 18636 26230 18642
rect 26256 18636 26259 18662
rect 22163 18606 22169 18623
rect 22186 18606 22192 18623
rect 22163 18603 22192 18606
rect 22211 18621 22248 18624
rect 22211 18604 22217 18621
rect 22234 18608 22248 18621
rect 22262 18623 22291 18626
rect 22234 18604 22240 18608
rect 22116 18602 22119 18603
rect 22211 18601 22240 18604
rect 22262 18606 22268 18623
rect 22285 18622 22291 18623
rect 22317 18622 22320 18628
rect 22285 18608 22320 18622
rect 22285 18606 22291 18608
rect 22262 18603 22291 18606
rect 22317 18602 22320 18608
rect 22346 18602 22349 18628
rect 21406 18574 21972 18588
rect 21306 18555 21335 18558
rect 21306 18538 21312 18555
rect 21329 18538 21335 18555
rect 21306 18535 21335 18538
rect 21351 18534 21354 18560
rect 21380 18534 21383 18560
rect 21958 18558 21972 18574
rect 23145 18568 23148 18594
rect 23174 18588 23177 18594
rect 24120 18588 24134 18636
rect 24157 18602 24160 18628
rect 24186 18622 24189 18628
rect 24250 18623 24279 18626
rect 24250 18622 24256 18623
rect 24186 18608 24256 18622
rect 24186 18602 24189 18608
rect 24250 18606 24256 18608
rect 24273 18606 24279 18623
rect 26090 18623 26119 18626
rect 24250 18603 24279 18606
rect 24488 18608 25537 18622
rect 24488 18594 24502 18608
rect 24479 18592 24482 18594
rect 24410 18589 24439 18592
rect 24410 18588 24416 18589
rect 23174 18574 24416 18588
rect 23174 18568 23177 18574
rect 24410 18572 24416 18574
rect 24433 18572 24439 18589
rect 24410 18569 24439 18572
rect 24461 18589 24482 18592
rect 24461 18572 24467 18589
rect 24461 18569 24482 18572
rect 24479 18568 24482 18569
rect 24508 18568 24511 18594
rect 21950 18555 21979 18558
rect 21950 18538 21956 18555
rect 21973 18538 21979 18555
rect 25523 18554 25537 18608
rect 26090 18606 26096 18623
rect 26113 18622 26119 18623
rect 26687 18622 26690 18628
rect 26113 18608 26690 18622
rect 26113 18606 26119 18608
rect 26090 18603 26119 18606
rect 26687 18602 26690 18608
rect 26716 18602 26719 18628
rect 27478 18626 27492 18676
rect 27975 18636 27978 18662
rect 28004 18636 28007 18662
rect 27470 18623 27499 18626
rect 27470 18606 27476 18623
rect 27493 18606 27499 18623
rect 27470 18603 27499 18606
rect 27561 18602 27564 18628
rect 27590 18626 27593 18628
rect 28297 18627 28300 18628
rect 28139 18626 28300 18627
rect 27590 18622 27594 18626
rect 28131 18623 28300 18626
rect 27590 18608 27612 18622
rect 27590 18603 27594 18608
rect 28131 18606 28137 18623
rect 28154 18613 28300 18623
rect 28154 18606 28160 18613
rect 28131 18603 28160 18606
rect 27590 18602 27593 18603
rect 28297 18602 28300 18613
rect 28326 18602 28329 18628
rect 26227 18568 26230 18594
rect 26256 18568 26259 18594
rect 26273 18568 26276 18594
rect 26302 18568 26305 18594
rect 27377 18568 27380 18594
rect 27406 18568 27409 18594
rect 27515 18568 27518 18594
rect 27544 18568 27547 18594
rect 28183 18589 28212 18592
rect 28183 18572 28189 18589
rect 28206 18588 28212 18589
rect 28251 18588 28254 18594
rect 28206 18574 28254 18588
rect 28206 18572 28212 18574
rect 28183 18569 28212 18572
rect 28251 18568 28254 18574
rect 28280 18568 28283 18594
rect 26457 18554 26460 18560
rect 25523 18540 26460 18554
rect 21950 18535 21979 18538
rect 26457 18534 26460 18540
rect 26486 18534 26489 18560
rect 28435 18534 28438 18560
rect 28464 18554 28467 18560
rect 29011 18555 29040 18558
rect 29011 18554 29017 18555
rect 28464 18540 29017 18554
rect 28464 18534 28467 18540
rect 29011 18538 29017 18540
rect 29034 18538 29040 18555
rect 29011 18535 29040 18538
rect 3036 18472 29992 18520
rect 4355 18453 4384 18456
rect 4355 18436 4361 18453
rect 4378 18452 4384 18453
rect 4791 18452 4794 18458
rect 4378 18438 4794 18452
rect 4378 18436 4384 18438
rect 4355 18433 4384 18436
rect 4791 18432 4794 18438
rect 4820 18432 4823 18458
rect 4837 18432 4840 18458
rect 4866 18452 4869 18458
rect 6033 18452 6036 18458
rect 4866 18438 6036 18452
rect 4866 18432 4869 18438
rect 6033 18432 6036 18438
rect 6062 18452 6065 18458
rect 6218 18453 6247 18456
rect 6218 18452 6224 18453
rect 6062 18438 6224 18452
rect 6062 18432 6065 18438
rect 6218 18436 6224 18438
rect 6241 18436 6247 18453
rect 6218 18433 6247 18436
rect 6263 18432 6266 18458
rect 6292 18432 6295 18458
rect 9529 18432 9532 18458
rect 9558 18452 9561 18458
rect 9558 18438 9667 18452
rect 9558 18432 9561 18438
rect 3549 18422 3552 18424
rect 3531 18419 3552 18422
rect 3531 18402 3537 18419
rect 3531 18399 3552 18402
rect 3549 18398 3552 18399
rect 3578 18398 3581 18424
rect 6889 18419 6918 18422
rect 6889 18402 6895 18419
rect 6912 18418 6918 18419
rect 9653 18418 9667 18438
rect 11001 18432 11004 18458
rect 11030 18456 11033 18458
rect 11030 18453 11054 18456
rect 11030 18436 11031 18453
rect 11048 18452 11054 18453
rect 11048 18438 11077 18452
rect 11048 18436 11054 18438
rect 11030 18433 11054 18436
rect 11030 18432 11033 18433
rect 11645 18432 11648 18458
rect 11674 18452 11677 18458
rect 12841 18452 12844 18458
rect 11674 18438 12844 18452
rect 11674 18432 11677 18438
rect 12841 18432 12844 18438
rect 12870 18432 12873 18458
rect 13991 18432 13994 18458
rect 14020 18452 14023 18458
rect 14451 18452 14454 18458
rect 14020 18438 14454 18452
rect 14020 18432 14023 18438
rect 14451 18432 14454 18438
rect 14480 18432 14483 18458
rect 15785 18432 15788 18458
rect 15814 18452 15817 18458
rect 16522 18453 16551 18456
rect 16522 18452 16528 18453
rect 15814 18438 16528 18452
rect 15814 18432 15817 18438
rect 16522 18436 16528 18438
rect 16545 18436 16551 18453
rect 16522 18433 16551 18436
rect 17165 18432 17168 18458
rect 17194 18432 17197 18458
rect 19351 18453 19380 18456
rect 19351 18436 19357 18453
rect 19374 18452 19380 18453
rect 20661 18452 20664 18458
rect 19374 18438 20664 18452
rect 19374 18436 19380 18438
rect 19351 18433 19380 18436
rect 20661 18432 20664 18438
rect 20690 18432 20693 18458
rect 21789 18453 21818 18456
rect 21789 18436 21795 18453
rect 21812 18452 21818 18453
rect 21949 18452 21952 18458
rect 21812 18438 21952 18452
rect 21812 18436 21818 18438
rect 21789 18433 21818 18436
rect 21949 18432 21952 18438
rect 21978 18432 21981 18458
rect 24043 18453 24072 18456
rect 24043 18436 24049 18453
rect 24066 18452 24072 18453
rect 24066 18438 24456 18452
rect 24066 18436 24072 18438
rect 24043 18433 24072 18436
rect 10219 18422 10222 18424
rect 10201 18419 10222 18422
rect 6912 18404 7022 18418
rect 9653 18404 9736 18418
rect 6912 18402 6918 18404
rect 6889 18399 6918 18402
rect 7008 18390 7022 18404
rect 3135 18364 3138 18390
rect 3164 18384 3167 18390
rect 3320 18385 3349 18388
rect 3320 18384 3326 18385
rect 3164 18370 3326 18384
rect 3164 18364 3167 18370
rect 3320 18368 3326 18370
rect 3343 18368 3349 18385
rect 3320 18365 3349 18368
rect 3481 18385 3510 18388
rect 3481 18368 3487 18385
rect 3504 18384 3510 18385
rect 3595 18384 3598 18390
rect 3504 18370 3598 18384
rect 3504 18368 3510 18370
rect 3481 18365 3510 18368
rect 3595 18364 3598 18370
rect 3624 18364 3627 18390
rect 5573 18364 5576 18390
rect 5602 18384 5605 18390
rect 6171 18384 6174 18390
rect 5602 18370 6174 18384
rect 5602 18364 5605 18370
rect 6171 18364 6174 18370
rect 6200 18384 6203 18390
rect 6839 18385 6868 18388
rect 6839 18384 6845 18385
rect 6200 18370 6845 18384
rect 6200 18364 6203 18370
rect 6839 18368 6845 18370
rect 6862 18384 6868 18385
rect 6953 18384 6956 18390
rect 6862 18370 6956 18384
rect 6862 18368 6868 18370
rect 6839 18365 6868 18368
rect 6953 18364 6956 18370
rect 6982 18364 6985 18390
rect 6999 18364 7002 18390
rect 7028 18384 7031 18390
rect 7091 18384 7094 18390
rect 7028 18370 7094 18384
rect 7028 18364 7031 18370
rect 7091 18364 7094 18370
rect 7120 18364 7123 18390
rect 9299 18364 9302 18390
rect 9328 18384 9331 18390
rect 9346 18385 9375 18388
rect 9346 18384 9352 18385
rect 9328 18370 9352 18384
rect 9328 18364 9331 18370
rect 9346 18368 9352 18370
rect 9369 18368 9375 18385
rect 9346 18365 9375 18368
rect 9391 18364 9394 18390
rect 9420 18388 9423 18390
rect 9420 18385 9432 18388
rect 9426 18368 9432 18385
rect 9420 18365 9432 18368
rect 9420 18364 9423 18365
rect 9483 18364 9486 18390
rect 9512 18388 9515 18390
rect 9512 18385 9526 18388
rect 9520 18368 9526 18385
rect 9544 18374 9547 18400
rect 9573 18374 9576 18400
rect 9607 18385 9636 18388
rect 9512 18365 9526 18368
rect 9607 18368 9613 18385
rect 9630 18384 9636 18385
rect 9658 18385 9687 18388
rect 9630 18368 9644 18384
rect 9607 18365 9644 18368
rect 9658 18368 9664 18385
rect 9681 18368 9687 18385
rect 9722 18384 9736 18404
rect 10201 18402 10207 18419
rect 10201 18399 10222 18402
rect 10219 18398 10222 18399
rect 10248 18398 10251 18424
rect 12795 18398 12798 18424
rect 12824 18418 12827 18424
rect 13003 18419 13032 18422
rect 13003 18418 13009 18419
rect 12824 18404 13009 18418
rect 12824 18398 12827 18404
rect 13003 18402 13009 18404
rect 13026 18402 13032 18419
rect 13003 18399 13032 18402
rect 15049 18398 15052 18424
rect 15078 18418 15081 18424
rect 15348 18419 15377 18422
rect 15348 18418 15354 18419
rect 15078 18404 15354 18418
rect 15078 18398 15081 18404
rect 15348 18402 15354 18404
rect 15371 18402 15377 18419
rect 15348 18399 15377 18402
rect 16223 18419 16252 18422
rect 16223 18402 16229 18419
rect 16246 18418 16252 18419
rect 17074 18419 17103 18422
rect 16246 18404 16590 18418
rect 16246 18402 16252 18404
rect 16223 18399 16252 18402
rect 10145 18385 10174 18388
rect 10145 18384 10151 18385
rect 9722 18370 10151 18384
rect 9658 18365 9687 18368
rect 10145 18368 10151 18370
rect 10168 18384 10174 18385
rect 10311 18384 10314 18390
rect 10168 18370 10314 18384
rect 10168 18368 10174 18370
rect 10145 18365 10174 18368
rect 9512 18364 9515 18365
rect 5389 18330 5392 18356
rect 5418 18350 5421 18356
rect 6310 18351 6339 18354
rect 6310 18350 6316 18351
rect 5418 18336 6316 18350
rect 5418 18330 5421 18336
rect 6310 18334 6316 18336
rect 6333 18334 6339 18351
rect 6310 18331 6339 18334
rect 6678 18351 6707 18354
rect 6678 18334 6684 18351
rect 6701 18334 6707 18351
rect 6678 18331 6707 18334
rect 5297 18262 5300 18288
rect 5326 18282 5329 18288
rect 6034 18283 6063 18286
rect 6034 18282 6040 18283
rect 5326 18268 6040 18282
rect 5326 18262 5329 18268
rect 6034 18266 6040 18268
rect 6057 18266 6063 18283
rect 6686 18282 6700 18331
rect 9346 18317 9375 18320
rect 9346 18300 9352 18317
rect 9369 18316 9375 18317
rect 9437 18316 9440 18322
rect 9369 18302 9440 18316
rect 9369 18300 9375 18302
rect 9346 18297 9375 18300
rect 9437 18296 9440 18302
rect 9466 18296 9469 18322
rect 9483 18296 9486 18322
rect 9512 18316 9515 18322
rect 9630 18316 9644 18365
rect 9512 18302 9644 18316
rect 9512 18296 9515 18302
rect 6953 18282 6956 18288
rect 6686 18268 6956 18282
rect 6034 18263 6063 18266
rect 6953 18262 6956 18268
rect 6982 18282 6985 18288
rect 7275 18282 7278 18288
rect 6982 18268 7278 18282
rect 6982 18262 6985 18268
rect 7275 18262 7278 18268
rect 7304 18262 7307 18288
rect 7505 18262 7508 18288
rect 7534 18282 7537 18288
rect 7713 18283 7742 18286
rect 7713 18282 7719 18283
rect 7534 18268 7719 18282
rect 7534 18262 7537 18268
rect 7713 18266 7719 18268
rect 7736 18266 7742 18283
rect 7713 18263 7742 18266
rect 9207 18262 9210 18288
rect 9236 18282 9239 18288
rect 9666 18282 9680 18365
rect 10311 18364 10314 18370
rect 10340 18364 10343 18390
rect 12957 18385 12986 18388
rect 12957 18368 12963 18385
rect 12980 18384 12986 18385
rect 13071 18384 13074 18390
rect 12980 18370 13074 18384
rect 12980 18368 12986 18370
rect 12957 18365 12986 18368
rect 13071 18364 13074 18370
rect 13100 18364 13103 18390
rect 13669 18364 13672 18390
rect 13698 18384 13701 18390
rect 15233 18384 15236 18390
rect 13698 18370 15236 18384
rect 13698 18364 13701 18370
rect 15233 18364 15236 18370
rect 15262 18364 15265 18390
rect 15387 18385 15416 18388
rect 15387 18368 15393 18385
rect 15410 18384 15416 18385
rect 15509 18384 15512 18390
rect 15410 18370 15512 18384
rect 15410 18368 15416 18370
rect 15387 18365 15416 18368
rect 15509 18364 15512 18370
rect 15538 18364 15541 18390
rect 15739 18364 15742 18390
rect 15768 18384 15771 18390
rect 16476 18385 16505 18388
rect 15768 18370 16452 18384
rect 15768 18364 15771 18370
rect 9990 18351 10019 18354
rect 9990 18334 9996 18351
rect 10013 18334 10019 18351
rect 9990 18331 10019 18334
rect 9236 18268 9680 18282
rect 9998 18282 10012 18331
rect 12749 18330 12752 18356
rect 12778 18350 12781 18356
rect 12796 18351 12825 18354
rect 12796 18350 12802 18351
rect 12778 18336 12802 18350
rect 12778 18330 12781 18336
rect 12796 18334 12802 18336
rect 12819 18334 12825 18351
rect 12796 18331 12825 18334
rect 14451 18330 14454 18356
rect 14480 18350 14483 18356
rect 15187 18350 15190 18356
rect 14480 18336 15190 18350
rect 14480 18330 14483 18336
rect 15187 18330 15190 18336
rect 15216 18330 15219 18356
rect 16438 18350 16452 18370
rect 16476 18368 16482 18385
rect 16499 18384 16505 18385
rect 16521 18384 16524 18390
rect 16499 18370 16524 18384
rect 16499 18368 16505 18370
rect 16476 18365 16505 18368
rect 16521 18364 16524 18370
rect 16550 18364 16553 18390
rect 16576 18388 16590 18404
rect 17074 18402 17080 18419
rect 17097 18418 17103 18419
rect 17174 18418 17188 18432
rect 17097 18404 17188 18418
rect 18527 18419 18556 18422
rect 17097 18402 17103 18404
rect 17074 18399 17103 18402
rect 18527 18402 18533 18419
rect 18550 18402 18556 18419
rect 18527 18399 18556 18402
rect 16568 18385 16597 18388
rect 16568 18368 16574 18385
rect 16591 18368 16597 18385
rect 16568 18365 16597 18368
rect 17119 18364 17122 18390
rect 17148 18384 17151 18390
rect 17166 18385 17195 18388
rect 17166 18384 17172 18385
rect 17148 18370 17172 18384
rect 17148 18364 17151 18370
rect 17166 18368 17172 18370
rect 17189 18368 17195 18385
rect 17166 18365 17195 18368
rect 17211 18364 17214 18390
rect 17240 18364 17243 18390
rect 17257 18364 17260 18390
rect 17286 18388 17289 18390
rect 17286 18384 17290 18388
rect 17286 18370 17308 18384
rect 17286 18365 17290 18370
rect 17286 18364 17289 18365
rect 17947 18364 17950 18390
rect 17976 18384 17979 18390
rect 18453 18384 18456 18390
rect 18482 18388 18485 18390
rect 18482 18385 18500 18388
rect 17976 18370 18456 18384
rect 17976 18364 17979 18370
rect 18453 18364 18456 18370
rect 18494 18368 18500 18385
rect 18534 18384 18548 18399
rect 23053 18398 23056 18424
rect 23082 18418 23085 18424
rect 23215 18419 23244 18422
rect 23215 18418 23221 18419
rect 23082 18404 23221 18418
rect 23082 18398 23085 18404
rect 23215 18402 23221 18404
rect 23238 18402 23244 18419
rect 23215 18399 23244 18402
rect 24295 18398 24298 18424
rect 24324 18398 24327 18424
rect 24442 18422 24456 18438
rect 27515 18432 27518 18458
rect 27544 18452 27547 18458
rect 28435 18452 28438 18458
rect 27544 18438 28438 18452
rect 27544 18432 27547 18438
rect 28435 18432 28438 18438
rect 28464 18432 28467 18458
rect 29425 18453 29454 18456
rect 29425 18436 29431 18453
rect 29448 18452 29454 18453
rect 29631 18452 29634 18458
rect 29448 18438 29634 18452
rect 29448 18436 29454 18438
rect 29425 18433 29454 18436
rect 29631 18432 29634 18438
rect 29660 18432 29663 18458
rect 24434 18419 24463 18422
rect 24434 18402 24440 18419
rect 24457 18402 24463 18419
rect 24434 18399 24463 18402
rect 28343 18398 28346 18424
rect 28372 18418 28375 18424
rect 28619 18422 28622 18424
rect 28550 18419 28579 18422
rect 28550 18418 28556 18419
rect 28372 18404 28556 18418
rect 28372 18398 28375 18404
rect 28550 18402 28556 18404
rect 28573 18402 28579 18419
rect 28550 18399 28579 18402
rect 28601 18419 28622 18422
rect 28601 18402 28607 18419
rect 28601 18399 28622 18402
rect 28619 18398 28622 18399
rect 28648 18398 28651 18424
rect 18913 18384 18916 18390
rect 18534 18370 18916 18384
rect 18482 18365 18500 18368
rect 18482 18364 18485 18365
rect 18913 18364 18916 18370
rect 18942 18364 18945 18390
rect 20661 18364 20664 18390
rect 20690 18384 20693 18390
rect 20909 18385 20938 18388
rect 20909 18384 20915 18385
rect 20690 18370 20915 18384
rect 20690 18364 20693 18370
rect 20909 18368 20915 18370
rect 20932 18368 20938 18385
rect 20909 18365 20938 18368
rect 20953 18385 20982 18388
rect 20953 18368 20959 18385
rect 20976 18384 20982 18385
rect 21305 18384 21308 18390
rect 20976 18370 21308 18384
rect 20976 18368 20982 18370
rect 20953 18365 20982 18368
rect 21305 18364 21308 18370
rect 21334 18384 21337 18390
rect 21627 18384 21630 18390
rect 21334 18370 21630 18384
rect 21334 18364 21337 18370
rect 21627 18364 21630 18370
rect 21656 18364 21659 18390
rect 22777 18364 22780 18390
rect 22806 18384 22809 18390
rect 23145 18384 23148 18390
rect 23174 18388 23177 18390
rect 23174 18385 23192 18388
rect 22806 18370 23148 18384
rect 22806 18364 22809 18370
rect 23145 18364 23148 18370
rect 23186 18368 23192 18385
rect 23174 18365 23192 18368
rect 23174 18364 23177 18365
rect 24387 18364 24390 18390
rect 24416 18364 24419 18390
rect 24479 18364 24482 18390
rect 24508 18388 24511 18390
rect 24508 18384 24512 18388
rect 27561 18384 27564 18390
rect 24508 18370 27564 18384
rect 24508 18365 24512 18370
rect 24508 18364 24511 18365
rect 27561 18364 27564 18370
rect 27590 18384 27593 18390
rect 29769 18384 29772 18390
rect 27590 18370 29772 18384
rect 27590 18364 27593 18370
rect 29769 18364 29772 18370
rect 29798 18364 29801 18390
rect 17074 18351 17103 18354
rect 17074 18350 17080 18351
rect 16438 18336 17080 18350
rect 17074 18334 17080 18336
rect 17097 18334 17103 18351
rect 17074 18331 17103 18334
rect 18316 18351 18345 18354
rect 18316 18334 18322 18351
rect 18339 18334 18345 18351
rect 18316 18331 18345 18334
rect 20754 18351 20783 18354
rect 20754 18334 20760 18351
rect 20777 18334 20783 18351
rect 20754 18331 20783 18334
rect 10173 18282 10176 18288
rect 9998 18268 10176 18282
rect 9236 18262 9239 18268
rect 10173 18262 10176 18268
rect 10202 18262 10205 18288
rect 13831 18283 13860 18286
rect 13831 18266 13837 18283
rect 13854 18282 13860 18283
rect 14681 18282 14684 18288
rect 13854 18268 14684 18282
rect 13854 18266 13860 18268
rect 13831 18263 13860 18266
rect 14681 18262 14684 18268
rect 14710 18262 14713 18288
rect 18324 18282 18338 18331
rect 19235 18282 19238 18288
rect 18324 18268 19238 18282
rect 19235 18262 19238 18268
rect 19264 18262 19267 18288
rect 20762 18282 20776 18331
rect 22961 18330 22964 18356
rect 22990 18350 22993 18356
rect 23008 18351 23037 18354
rect 23008 18350 23014 18351
rect 22990 18336 23014 18350
rect 22990 18330 22993 18336
rect 23008 18334 23014 18336
rect 23031 18334 23037 18351
rect 23008 18331 23037 18334
rect 21075 18282 21078 18288
rect 20762 18268 21078 18282
rect 21075 18262 21078 18268
rect 21104 18262 21107 18288
rect 23016 18282 23030 18331
rect 24341 18330 24344 18356
rect 24370 18330 24373 18356
rect 24396 18350 24410 18364
rect 24396 18336 24502 18350
rect 24488 18322 24502 18336
rect 27975 18330 27978 18356
rect 28004 18350 28007 18356
rect 28390 18351 28419 18354
rect 28390 18350 28396 18351
rect 28004 18336 28396 18350
rect 28004 18330 28007 18336
rect 28390 18334 28396 18336
rect 28413 18334 28419 18351
rect 28390 18331 28419 18334
rect 24479 18296 24482 18322
rect 24508 18296 24511 18322
rect 23145 18282 23148 18288
rect 23016 18268 23148 18282
rect 23145 18262 23148 18268
rect 23174 18282 23177 18288
rect 24157 18282 24160 18288
rect 23174 18268 24160 18282
rect 23174 18262 23177 18268
rect 24157 18262 24160 18268
rect 24186 18262 24189 18288
rect 3036 18200 29992 18248
rect 3595 18180 3598 18186
rect 3144 18166 3598 18180
rect 3144 18112 3158 18166
rect 3595 18160 3598 18166
rect 3624 18160 3627 18186
rect 4171 18181 4200 18184
rect 4171 18164 4177 18181
rect 4194 18180 4200 18181
rect 4653 18180 4656 18186
rect 4194 18166 4656 18180
rect 4194 18164 4200 18166
rect 4171 18161 4200 18164
rect 4653 18160 4656 18166
rect 4682 18160 4685 18186
rect 5665 18180 5668 18186
rect 5214 18166 5668 18180
rect 5160 18113 5189 18116
rect 3144 18098 3204 18112
rect 3135 18058 3138 18084
rect 3164 18058 3167 18084
rect 3190 18078 3204 18098
rect 5160 18096 5166 18113
rect 5183 18112 5189 18113
rect 5214 18112 5228 18166
rect 5665 18160 5668 18166
rect 5694 18160 5697 18186
rect 6033 18160 6036 18186
rect 6062 18160 6065 18186
rect 6907 18160 6910 18186
rect 6936 18180 6939 18186
rect 7414 18181 7443 18184
rect 7414 18180 7420 18181
rect 6936 18166 7420 18180
rect 6936 18160 6939 18166
rect 7414 18164 7420 18166
rect 7437 18164 7443 18181
rect 9115 18180 9118 18186
rect 7414 18161 7443 18164
rect 8434 18166 9118 18180
rect 6769 18126 6772 18152
rect 6798 18146 6801 18152
rect 8434 18146 8448 18166
rect 9115 18160 9118 18166
rect 9144 18180 9147 18186
rect 9483 18184 9486 18186
rect 9461 18181 9486 18184
rect 9144 18166 9276 18180
rect 9144 18160 9147 18166
rect 6798 18132 8448 18146
rect 9262 18146 9276 18166
rect 9461 18164 9467 18181
rect 9484 18164 9486 18181
rect 9461 18161 9486 18164
rect 9483 18160 9486 18161
rect 9512 18160 9515 18186
rect 10771 18180 10774 18186
rect 10182 18166 10774 18180
rect 10182 18146 10196 18166
rect 10771 18160 10774 18166
rect 10800 18160 10803 18186
rect 10863 18160 10866 18186
rect 10892 18180 10895 18186
rect 11209 18181 11238 18184
rect 11209 18180 11215 18181
rect 10892 18166 11215 18180
rect 10892 18160 10895 18166
rect 11209 18164 11215 18166
rect 11232 18164 11238 18181
rect 13853 18180 13856 18186
rect 11209 18161 11238 18164
rect 13402 18166 13856 18180
rect 9262 18132 10196 18146
rect 6798 18126 6801 18132
rect 5183 18098 5228 18112
rect 5183 18096 5189 18098
rect 5160 18093 5189 18096
rect 5297 18092 5300 18118
rect 5326 18092 5329 18118
rect 7551 18092 7554 18118
rect 7580 18112 7583 18118
rect 7580 18098 7942 18112
rect 7580 18092 7583 18098
rect 3291 18079 3320 18082
rect 3291 18078 3297 18079
rect 3190 18064 3297 18078
rect 3291 18062 3297 18064
rect 3314 18062 3320 18079
rect 3733 18078 3736 18084
rect 3291 18059 3320 18062
rect 3354 18064 3736 18078
rect 3354 18048 3368 18064
rect 3733 18058 3736 18064
rect 3762 18058 3765 18084
rect 6677 18058 6680 18084
rect 6706 18058 6709 18084
rect 6723 18058 6726 18084
rect 6752 18078 6755 18084
rect 6861 18078 6864 18084
rect 6752 18064 6864 18078
rect 6752 18058 6755 18064
rect 6861 18058 6864 18064
rect 6890 18058 6893 18084
rect 7414 18079 7443 18082
rect 7414 18078 7420 18079
rect 6962 18064 7420 18078
rect 3347 18045 3376 18048
rect 3347 18028 3353 18045
rect 3370 18028 3376 18045
rect 3347 18025 3376 18028
rect 5573 18024 5576 18050
rect 5602 18024 5605 18050
rect 5987 18044 5990 18050
rect 5911 18030 5990 18044
rect 5987 18024 5990 18030
rect 6016 18024 6019 18050
rect 6769 18024 6772 18050
rect 6798 18024 6801 18050
rect 6815 18024 6818 18050
rect 6844 18024 6847 18050
rect 6962 18014 6976 18064
rect 7414 18062 7420 18064
rect 7437 18062 7443 18079
rect 7414 18059 7443 18062
rect 7460 18079 7489 18082
rect 7460 18062 7466 18079
rect 7483 18078 7489 18079
rect 7505 18078 7508 18084
rect 7483 18064 7508 18078
rect 7483 18062 7489 18064
rect 7460 18059 7489 18062
rect 7505 18058 7508 18064
rect 7534 18058 7537 18084
rect 7643 18058 7646 18084
rect 7672 18058 7675 18084
rect 7552 18045 7581 18048
rect 7552 18028 7558 18045
rect 7575 18028 7581 18045
rect 7552 18025 7581 18028
rect 6954 18011 6983 18014
rect 6954 17994 6960 18011
rect 6977 17994 6983 18011
rect 7560 18010 7574 18025
rect 7597 18024 7600 18050
rect 7626 18024 7629 18050
rect 7928 18044 7942 18098
rect 8287 18058 8290 18084
rect 8316 18078 8319 18084
rect 8425 18078 8428 18084
rect 8316 18064 8428 18078
rect 8316 18058 8319 18064
rect 8425 18058 8428 18064
rect 8454 18058 8457 18084
rect 8563 18058 8566 18084
rect 8592 18082 8595 18084
rect 8592 18079 8610 18082
rect 8604 18062 8610 18079
rect 8592 18059 8610 18062
rect 8592 18058 8595 18059
rect 10173 18058 10176 18084
rect 10202 18058 10205 18084
rect 10311 18058 10314 18084
rect 10340 18082 10343 18084
rect 10340 18079 10358 18082
rect 10352 18062 10358 18079
rect 10340 18059 10358 18062
rect 10340 18058 10343 18059
rect 12749 18058 12752 18084
rect 12778 18078 12781 18084
rect 13402 18082 13416 18166
rect 13853 18160 13856 18166
rect 13882 18180 13885 18186
rect 14451 18180 14454 18186
rect 13882 18166 14454 18180
rect 13882 18160 13885 18166
rect 14451 18160 14454 18166
rect 14480 18160 14483 18186
rect 14681 18160 14684 18186
rect 14710 18180 14713 18186
rect 14710 18166 14965 18180
rect 14710 18160 14713 18166
rect 14865 18126 14868 18152
rect 14894 18146 14897 18152
rect 14894 18126 14903 18146
rect 14429 18113 14458 18116
rect 14429 18096 14435 18113
rect 14452 18112 14458 18113
rect 14452 18098 14842 18112
rect 14452 18096 14458 18098
rect 14429 18093 14458 18096
rect 13394 18079 13423 18082
rect 13394 18078 13400 18079
rect 12778 18064 13400 18078
rect 12778 18058 12781 18064
rect 13394 18062 13400 18064
rect 13417 18062 13423 18079
rect 13555 18079 13584 18082
rect 13555 18078 13561 18079
rect 13394 18059 13423 18062
rect 13448 18064 13561 18078
rect 8333 18044 8336 18050
rect 7928 18030 8336 18044
rect 8333 18024 8336 18030
rect 8362 18044 8365 18050
rect 10403 18048 10406 18050
rect 8625 18045 8654 18048
rect 8625 18044 8631 18045
rect 8362 18030 8631 18044
rect 8362 18024 8365 18030
rect 8625 18028 8631 18030
rect 8648 18028 8654 18045
rect 8625 18025 8654 18028
rect 10385 18045 10406 18048
rect 10385 18028 10391 18045
rect 10385 18025 10406 18028
rect 10403 18024 10406 18025
rect 10432 18024 10435 18050
rect 12933 18024 12936 18050
rect 12962 18044 12965 18050
rect 13071 18044 13074 18050
rect 12962 18030 13074 18044
rect 12962 18024 12965 18030
rect 13071 18024 13074 18030
rect 13100 18044 13103 18050
rect 13448 18044 13462 18064
rect 13555 18062 13561 18064
rect 13578 18078 13584 18079
rect 13945 18078 13948 18084
rect 13578 18064 13948 18078
rect 13578 18062 13584 18064
rect 13555 18059 13584 18062
rect 13945 18058 13948 18064
rect 13974 18058 13977 18084
rect 14681 18058 14684 18084
rect 14710 18058 14713 18084
rect 14773 18082 14776 18084
rect 14759 18079 14776 18082
rect 14759 18062 14765 18079
rect 14759 18059 14776 18062
rect 14773 18058 14776 18059
rect 14802 18058 14805 18084
rect 14828 18082 14842 18098
rect 14889 18082 14903 18126
rect 14951 18088 14965 18166
rect 17211 18160 17214 18186
rect 17240 18184 17243 18186
rect 17240 18181 17264 18184
rect 17240 18164 17241 18181
rect 17258 18164 17264 18181
rect 17240 18161 17264 18164
rect 17240 18160 17243 18161
rect 20523 18160 20526 18186
rect 20552 18180 20555 18186
rect 20552 18166 20707 18180
rect 20552 18160 20555 18166
rect 15187 18092 15190 18118
rect 15216 18112 15219 18118
rect 20693 18112 20707 18166
rect 21121 18160 21124 18186
rect 21150 18180 21153 18186
rect 21351 18180 21354 18186
rect 21150 18166 21354 18180
rect 21150 18160 21153 18166
rect 21351 18160 21354 18166
rect 21380 18160 21383 18186
rect 21443 18160 21446 18186
rect 21472 18180 21475 18186
rect 21581 18180 21584 18186
rect 21472 18166 21584 18180
rect 21472 18160 21475 18166
rect 21581 18160 21584 18166
rect 21610 18160 21613 18186
rect 22087 18160 22090 18186
rect 22116 18180 22119 18186
rect 22249 18181 22278 18184
rect 22249 18180 22255 18181
rect 22116 18166 22255 18180
rect 22116 18160 22119 18166
rect 22249 18164 22255 18166
rect 22272 18164 22278 18181
rect 22249 18161 22278 18164
rect 23053 18160 23056 18186
rect 23082 18180 23085 18186
rect 28297 18180 28300 18186
rect 23082 18166 28300 18180
rect 23082 18160 23085 18166
rect 28297 18160 28300 18166
rect 28326 18180 28329 18186
rect 28435 18180 28438 18186
rect 28326 18166 28438 18180
rect 28326 18160 28329 18166
rect 28435 18160 28438 18166
rect 28464 18160 28467 18186
rect 22317 18126 22320 18152
rect 22346 18146 22349 18152
rect 27101 18146 27104 18152
rect 22346 18132 27104 18146
rect 22346 18126 22349 18132
rect 27101 18126 27104 18132
rect 27130 18126 27133 18152
rect 15216 18098 15877 18112
rect 20693 18098 21282 18112
rect 15216 18092 15219 18098
rect 14943 18085 14972 18088
rect 14828 18079 14862 18082
rect 14828 18064 14839 18079
rect 14833 18062 14839 18064
rect 14856 18062 14862 18079
rect 14833 18059 14862 18062
rect 14881 18079 14910 18082
rect 14881 18062 14887 18079
rect 14904 18062 14910 18079
rect 14943 18068 14949 18085
rect 14966 18068 14972 18085
rect 15003 18082 15006 18084
rect 14943 18065 14972 18068
rect 14994 18079 15006 18082
rect 14881 18059 14910 18062
rect 14994 18062 15000 18079
rect 14994 18059 15006 18062
rect 15003 18058 15006 18059
rect 15032 18058 15035 18084
rect 15049 18058 15052 18084
rect 15078 18058 15081 18084
rect 15863 18078 15877 18098
rect 16153 18078 16156 18084
rect 15863 18064 16156 18078
rect 16153 18058 16156 18064
rect 16182 18078 16185 18084
rect 16200 18079 16229 18082
rect 16200 18078 16206 18079
rect 16182 18064 16206 18078
rect 16182 18058 16185 18064
rect 16200 18062 16206 18064
rect 16223 18078 16229 18079
rect 17717 18078 17720 18084
rect 16223 18064 17720 18078
rect 16223 18062 16229 18064
rect 16200 18059 16229 18062
rect 17717 18058 17720 18064
rect 17746 18058 17749 18084
rect 20661 18058 20664 18084
rect 20690 18078 20693 18084
rect 20690 18058 20707 18078
rect 21075 18058 21078 18084
rect 21104 18078 21107 18084
rect 21214 18079 21243 18082
rect 21214 18078 21220 18079
rect 21104 18064 21220 18078
rect 21104 18058 21107 18064
rect 21214 18062 21220 18064
rect 21237 18062 21243 18079
rect 21268 18078 21282 18098
rect 23237 18092 23240 18118
rect 23266 18112 23269 18118
rect 23421 18112 23424 18118
rect 23266 18098 23424 18112
rect 23266 18092 23269 18098
rect 23421 18092 23424 18098
rect 23450 18092 23453 18118
rect 21627 18078 21630 18084
rect 21268 18064 21630 18078
rect 21214 18059 21243 18062
rect 21627 18058 21630 18064
rect 21656 18058 21659 18084
rect 13623 18048 13626 18050
rect 13100 18030 13462 18044
rect 13605 18045 13626 18048
rect 13100 18024 13103 18030
rect 13605 18028 13611 18045
rect 13605 18025 13626 18028
rect 13623 18024 13626 18025
rect 13652 18024 13655 18050
rect 15058 18044 15072 18058
rect 16360 18045 16389 18048
rect 16360 18044 16366 18045
rect 15058 18030 16366 18044
rect 16360 18028 16366 18030
rect 16383 18028 16389 18045
rect 16360 18025 16389 18028
rect 16411 18045 16440 18048
rect 16411 18028 16417 18045
rect 16434 18044 16440 18045
rect 16475 18044 16478 18050
rect 16434 18030 16478 18044
rect 16434 18028 16440 18030
rect 16411 18025 16440 18028
rect 16475 18024 16478 18030
rect 16504 18024 16507 18050
rect 20693 18044 20707 18058
rect 21443 18048 21446 18050
rect 21374 18045 21403 18048
rect 21374 18044 21380 18045
rect 20693 18030 21380 18044
rect 21374 18028 21380 18030
rect 21397 18028 21403 18045
rect 21374 18025 21403 18028
rect 21425 18045 21446 18048
rect 21425 18028 21431 18045
rect 21425 18025 21446 18028
rect 21443 18024 21446 18025
rect 21472 18024 21475 18050
rect 7689 18010 7692 18016
rect 7560 17996 7692 18010
rect 6954 17991 6983 17994
rect 7689 17990 7692 17996
rect 7718 17990 7721 18016
rect 14912 18011 14941 18014
rect 14912 17994 14918 18011
rect 14935 18010 14941 18011
rect 15049 18010 15052 18016
rect 14935 17996 15052 18010
rect 14935 17994 14941 17996
rect 14912 17991 14941 17994
rect 15049 17990 15052 17996
rect 15078 17990 15081 18016
rect 19373 17990 19376 18016
rect 19402 18010 19405 18016
rect 20155 18010 20158 18016
rect 19402 17996 20158 18010
rect 19402 17990 19405 17996
rect 20155 17990 20158 17996
rect 20184 17990 20187 18016
rect 3036 17928 29992 17976
rect 13831 17909 13860 17912
rect 13831 17892 13837 17909
rect 13854 17908 13860 17909
rect 14681 17908 14684 17914
rect 13854 17894 14684 17908
rect 13854 17892 13860 17894
rect 13831 17889 13860 17892
rect 14681 17888 14684 17894
rect 14710 17888 14713 17914
rect 22111 17909 22140 17912
rect 22111 17892 22117 17909
rect 22134 17908 22140 17909
rect 22363 17908 22366 17914
rect 22134 17894 22366 17908
rect 22134 17892 22140 17894
rect 22111 17889 22140 17892
rect 22363 17888 22366 17894
rect 22392 17888 22395 17914
rect 24249 17888 24252 17914
rect 24278 17888 24281 17914
rect 5757 17854 5760 17880
rect 5786 17874 5789 17880
rect 6171 17874 6174 17880
rect 5786 17860 6174 17874
rect 5786 17854 5789 17860
rect 6171 17854 6174 17860
rect 6200 17874 6203 17880
rect 6838 17875 6867 17878
rect 6838 17874 6844 17875
rect 6200 17860 6844 17874
rect 6200 17854 6203 17860
rect 6838 17858 6844 17860
rect 6861 17858 6867 17875
rect 6838 17855 6867 17858
rect 6889 17875 6918 17878
rect 6889 17858 6895 17875
rect 6912 17874 6918 17875
rect 6912 17860 7022 17874
rect 6912 17858 6918 17860
rect 6889 17855 6918 17858
rect 7008 17846 7022 17860
rect 12427 17854 12430 17880
rect 12456 17874 12459 17880
rect 13007 17875 13036 17878
rect 13007 17874 13013 17875
rect 12456 17860 13013 17874
rect 12456 17854 12459 17860
rect 13007 17858 13013 17860
rect 13030 17874 13036 17875
rect 13071 17874 13074 17880
rect 13030 17860 13074 17874
rect 13030 17858 13036 17860
rect 13007 17855 13036 17858
rect 13071 17854 13074 17860
rect 13100 17854 13103 17880
rect 21287 17875 21316 17878
rect 21287 17858 21293 17875
rect 21310 17874 21316 17875
rect 21351 17874 21354 17880
rect 21310 17860 21354 17874
rect 21310 17858 21316 17860
rect 21287 17855 21316 17858
rect 21351 17854 21354 17860
rect 21380 17854 21383 17880
rect 22961 17878 22964 17880
rect 22943 17875 22964 17878
rect 22943 17858 22949 17875
rect 22943 17855 22964 17858
rect 22961 17854 22964 17855
rect 22990 17854 22993 17880
rect 26457 17878 26460 17880
rect 26439 17875 26460 17878
rect 26439 17858 26445 17875
rect 26439 17855 26460 17858
rect 26457 17854 26460 17855
rect 26486 17854 26489 17880
rect 6678 17841 6707 17844
rect 6678 17824 6684 17841
rect 6701 17840 6707 17841
rect 6953 17840 6956 17846
rect 6701 17826 6956 17840
rect 6701 17824 6707 17826
rect 6678 17821 6707 17824
rect 6953 17820 6956 17826
rect 6982 17820 6985 17846
rect 6999 17820 7002 17846
rect 7028 17820 7031 17846
rect 12749 17820 12752 17846
rect 12778 17840 12781 17846
rect 12796 17841 12825 17844
rect 12796 17840 12802 17841
rect 12778 17826 12802 17840
rect 12778 17820 12781 17826
rect 12796 17824 12802 17826
rect 12819 17824 12825 17841
rect 12796 17821 12825 17824
rect 12933 17820 12936 17846
rect 12962 17844 12965 17846
rect 12962 17841 12980 17844
rect 12974 17824 12980 17841
rect 12962 17821 12980 17824
rect 12962 17820 12965 17821
rect 18775 17820 18778 17846
rect 18804 17820 18807 17846
rect 18867 17820 18870 17846
rect 18896 17820 18899 17846
rect 20155 17820 20158 17846
rect 20184 17840 20187 17846
rect 20661 17840 20664 17846
rect 20184 17826 20664 17840
rect 20184 17820 20187 17826
rect 20661 17820 20664 17826
rect 20690 17840 20693 17846
rect 21237 17841 21266 17844
rect 21237 17840 21243 17841
rect 20690 17826 21243 17840
rect 20690 17820 20693 17826
rect 21237 17824 21243 17826
rect 21260 17840 21266 17841
rect 21489 17840 21492 17846
rect 21260 17826 21492 17840
rect 21260 17824 21266 17826
rect 21237 17821 21266 17824
rect 21489 17820 21492 17826
rect 21518 17820 21521 17846
rect 22777 17820 22780 17846
rect 22806 17840 22809 17846
rect 22887 17841 22916 17844
rect 22887 17840 22893 17841
rect 22806 17826 22893 17840
rect 22806 17820 22809 17826
rect 22887 17824 22893 17826
rect 22910 17824 22916 17841
rect 22887 17821 22916 17824
rect 23973 17820 23976 17846
rect 24002 17840 24005 17846
rect 24020 17841 24049 17844
rect 24020 17840 24026 17841
rect 24002 17826 24026 17840
rect 24002 17820 24005 17826
rect 24020 17824 24026 17826
rect 24043 17824 24049 17841
rect 24020 17821 24049 17824
rect 24065 17820 24068 17846
rect 24094 17844 24097 17846
rect 24094 17841 24106 17844
rect 24100 17824 24106 17841
rect 24171 17841 24200 17844
rect 24171 17840 24177 17841
rect 24094 17821 24106 17824
rect 24166 17824 24177 17840
rect 24194 17824 24200 17841
rect 24166 17821 24200 17824
rect 24233 17841 24262 17844
rect 24233 17824 24239 17841
rect 24256 17824 24262 17841
rect 24233 17821 24262 17824
rect 24281 17841 24310 17844
rect 24281 17824 24287 17841
rect 24304 17824 24310 17841
rect 24281 17821 24310 17824
rect 24332 17841 24361 17844
rect 24332 17824 24338 17841
rect 24355 17840 24361 17841
rect 26135 17840 26138 17846
rect 24355 17826 26138 17840
rect 24355 17824 24361 17826
rect 24332 17821 24361 17824
rect 24094 17820 24097 17821
rect 7597 17786 7600 17812
rect 7626 17806 7629 17812
rect 7713 17807 7742 17810
rect 7713 17806 7719 17807
rect 7626 17792 7719 17806
rect 7626 17786 7629 17792
rect 7713 17790 7719 17792
rect 7736 17790 7742 17807
rect 7713 17787 7742 17790
rect 21075 17786 21078 17812
rect 21104 17786 21107 17812
rect 22732 17807 22761 17810
rect 22732 17790 22738 17807
rect 22755 17790 22761 17807
rect 22732 17787 22761 17790
rect 23767 17807 23796 17810
rect 23767 17790 23773 17807
rect 23790 17806 23796 17807
rect 24166 17806 24180 17821
rect 23790 17792 24180 17806
rect 24241 17806 24255 17821
rect 24241 17792 24272 17806
rect 23790 17790 23796 17792
rect 23767 17787 23796 17790
rect 18822 17739 18851 17742
rect 18822 17722 18828 17739
rect 18845 17738 18851 17739
rect 19281 17738 19284 17744
rect 18845 17724 19284 17738
rect 18845 17722 18851 17724
rect 18822 17719 18851 17722
rect 19281 17718 19284 17724
rect 19310 17718 19313 17744
rect 21213 17718 21216 17744
rect 21242 17738 21245 17744
rect 21351 17738 21354 17744
rect 21242 17724 21354 17738
rect 21242 17718 21245 17724
rect 21351 17718 21354 17724
rect 21380 17718 21383 17744
rect 22455 17718 22458 17744
rect 22484 17738 22487 17744
rect 22740 17738 22754 17787
rect 23145 17738 23148 17744
rect 22484 17724 23148 17738
rect 22484 17718 22487 17724
rect 23145 17718 23148 17724
rect 23174 17718 23177 17744
rect 24258 17738 24272 17792
rect 24289 17778 24303 17821
rect 26135 17820 26138 17826
rect 26164 17820 26167 17846
rect 26365 17820 26368 17846
rect 26394 17844 26397 17846
rect 26394 17841 26412 17844
rect 26406 17824 26412 17841
rect 26394 17821 26412 17824
rect 26394 17820 26397 17821
rect 26181 17786 26184 17812
rect 26210 17806 26213 17812
rect 26228 17807 26257 17810
rect 26228 17806 26234 17807
rect 26210 17792 26234 17806
rect 26210 17786 26213 17792
rect 26228 17790 26234 17792
rect 26251 17790 26257 17807
rect 26228 17787 26257 17790
rect 27101 17786 27104 17812
rect 27130 17806 27133 17812
rect 27423 17806 27426 17812
rect 27130 17792 27426 17806
rect 27130 17786 27133 17792
rect 27423 17786 27426 17792
rect 27452 17786 27455 17812
rect 24289 17758 24298 17778
rect 24295 17752 24298 17758
rect 24324 17752 24327 17778
rect 29585 17772 29588 17778
rect 27041 17758 29588 17772
rect 25721 17738 25724 17744
rect 24258 17724 25724 17738
rect 25721 17718 25724 17724
rect 25750 17738 25753 17744
rect 27041 17738 27055 17758
rect 29585 17752 29588 17758
rect 29614 17752 29617 17778
rect 25750 17724 27055 17738
rect 25750 17718 25753 17724
rect 27101 17718 27104 17744
rect 27130 17738 27133 17744
rect 27263 17739 27292 17742
rect 27263 17738 27269 17739
rect 27130 17724 27269 17738
rect 27130 17718 27133 17724
rect 27263 17722 27269 17724
rect 27286 17722 27292 17739
rect 27263 17719 27292 17722
rect 3036 17656 29992 17704
rect 4654 17637 4683 17640
rect 4654 17620 4660 17637
rect 4677 17636 4683 17637
rect 4699 17636 4702 17642
rect 4677 17622 4702 17636
rect 4677 17620 4683 17622
rect 4654 17617 4683 17620
rect 4699 17616 4702 17622
rect 4728 17616 4731 17642
rect 6655 17637 6684 17640
rect 6655 17620 6661 17637
rect 6678 17636 6684 17637
rect 6815 17636 6818 17642
rect 6678 17622 6818 17636
rect 6678 17620 6684 17622
rect 6655 17617 6684 17620
rect 6815 17616 6818 17622
rect 6844 17616 6847 17642
rect 8425 17636 8428 17642
rect 8250 17622 8428 17636
rect 3135 17548 3138 17574
rect 3164 17548 3167 17574
rect 8250 17572 8264 17622
rect 8425 17616 8428 17622
rect 8454 17616 8457 17642
rect 9277 17637 9306 17640
rect 9277 17620 9283 17637
rect 9300 17636 9306 17637
rect 9391 17636 9394 17642
rect 9300 17622 9394 17636
rect 9300 17620 9306 17622
rect 9277 17617 9306 17620
rect 9391 17616 9394 17622
rect 9420 17616 9423 17642
rect 18775 17616 18778 17642
rect 18804 17616 18807 17642
rect 22915 17636 22918 17642
rect 20693 17622 22918 17636
rect 19005 17582 19008 17608
rect 19034 17602 19037 17608
rect 20109 17602 20112 17608
rect 19034 17588 20112 17602
rect 19034 17582 19037 17588
rect 20109 17582 20112 17588
rect 20138 17582 20141 17608
rect 8242 17569 8271 17572
rect 8242 17552 8248 17569
rect 8265 17552 8271 17569
rect 19143 17568 19146 17574
rect 8242 17549 8271 17552
rect 19045 17554 19146 17568
rect 3181 17514 3184 17540
rect 3210 17534 3213 17540
rect 3210 17520 3368 17534
rect 3210 17514 3213 17520
rect 3354 17504 3368 17520
rect 4745 17514 4748 17540
rect 4774 17514 4777 17540
rect 4856 17535 4885 17538
rect 4856 17518 4862 17535
rect 4879 17534 4885 17535
rect 5205 17534 5208 17540
rect 4879 17520 5208 17534
rect 4879 17518 4885 17520
rect 4856 17515 4885 17518
rect 5205 17514 5208 17520
rect 5234 17514 5237 17540
rect 5620 17535 5649 17538
rect 5620 17518 5626 17535
rect 5643 17534 5649 17535
rect 5665 17534 5668 17540
rect 5643 17520 5668 17534
rect 5643 17518 5649 17520
rect 5620 17515 5649 17518
rect 5665 17514 5668 17520
rect 5694 17514 5697 17540
rect 5757 17514 5760 17540
rect 5786 17538 5789 17540
rect 5786 17535 5804 17538
rect 5798 17518 5804 17535
rect 5786 17515 5804 17518
rect 8403 17535 8432 17538
rect 8403 17518 8409 17535
rect 8426 17534 8432 17535
rect 8563 17534 8566 17540
rect 8426 17520 8566 17534
rect 8426 17518 8432 17520
rect 8403 17515 8432 17518
rect 5786 17514 5789 17515
rect 8563 17514 8566 17520
rect 8592 17514 8595 17540
rect 18776 17535 18805 17538
rect 18776 17518 18782 17535
rect 18799 17518 18805 17535
rect 18776 17515 18805 17518
rect 3296 17501 3325 17504
rect 3296 17500 3302 17501
rect 3006 17486 3302 17500
rect 3006 17330 3020 17486
rect 3296 17484 3302 17486
rect 3319 17484 3325 17501
rect 3296 17481 3325 17484
rect 3347 17501 3376 17504
rect 3347 17484 3353 17501
rect 3370 17500 3376 17501
rect 3411 17500 3414 17506
rect 3370 17486 3414 17500
rect 3370 17484 3376 17486
rect 3347 17481 3376 17484
rect 3411 17480 3414 17486
rect 3440 17480 3443 17506
rect 4171 17501 4200 17504
rect 4171 17484 4177 17501
rect 4194 17500 4200 17501
rect 4654 17501 4683 17504
rect 4654 17500 4660 17501
rect 4194 17486 4660 17500
rect 4194 17484 4200 17486
rect 4171 17481 4200 17484
rect 4654 17484 4660 17486
rect 4677 17484 4683 17501
rect 4654 17481 4683 17484
rect 4791 17480 4794 17506
rect 4820 17480 4823 17506
rect 5849 17504 5852 17506
rect 5831 17501 5852 17504
rect 5831 17484 5837 17501
rect 5831 17481 5852 17484
rect 5849 17480 5852 17481
rect 5878 17480 5881 17506
rect 8471 17504 8474 17506
rect 8453 17501 8474 17504
rect 8453 17484 8459 17501
rect 8453 17481 8474 17484
rect 8471 17480 8474 17481
rect 8500 17480 8503 17506
rect 11185 17446 11188 17472
rect 11214 17466 11217 17472
rect 13899 17466 13902 17472
rect 11214 17452 13902 17466
rect 11214 17446 11217 17452
rect 13899 17446 13902 17452
rect 13928 17466 13931 17472
rect 14451 17466 14454 17472
rect 13928 17452 14454 17466
rect 13928 17446 13931 17452
rect 14451 17446 14454 17452
rect 14480 17466 14483 17472
rect 16199 17466 16202 17472
rect 14480 17452 16202 17466
rect 14480 17446 14483 17452
rect 16199 17446 16202 17452
rect 16228 17446 16231 17472
rect 18784 17466 18798 17515
rect 18821 17514 18824 17540
rect 18850 17538 18853 17540
rect 18850 17535 18862 17538
rect 18856 17518 18862 17535
rect 18850 17515 18862 17518
rect 18850 17514 18853 17515
rect 18913 17514 18916 17540
rect 18942 17538 18945 17540
rect 18942 17535 18956 17538
rect 19045 17536 19059 17554
rect 19143 17548 19146 17554
rect 19172 17548 19175 17574
rect 18950 17518 18956 17535
rect 19037 17533 19066 17536
rect 18942 17515 18956 17518
rect 18942 17514 18945 17515
rect 18988 17503 18991 17529
rect 19017 17503 19020 17529
rect 19037 17516 19043 17533
rect 19060 17516 19066 17533
rect 19037 17513 19066 17516
rect 19088 17535 19117 17538
rect 19088 17518 19094 17535
rect 19111 17534 19117 17535
rect 19925 17534 19928 17540
rect 19111 17520 19928 17534
rect 19111 17518 19117 17520
rect 19088 17515 19117 17518
rect 19925 17514 19928 17520
rect 19954 17534 19957 17540
rect 20693 17534 20707 17622
rect 22915 17616 22918 17622
rect 22944 17616 22947 17642
rect 23491 17637 23520 17640
rect 23491 17620 23497 17637
rect 23514 17636 23520 17637
rect 24065 17636 24068 17642
rect 23514 17622 24068 17636
rect 23514 17620 23520 17622
rect 23491 17617 23520 17620
rect 24065 17616 24068 17622
rect 24094 17616 24097 17642
rect 25768 17637 25797 17640
rect 24120 17622 25537 17636
rect 23973 17582 23976 17608
rect 24002 17602 24005 17608
rect 24120 17602 24134 17622
rect 24002 17588 24134 17602
rect 24002 17582 24005 17588
rect 21075 17548 21078 17574
rect 21104 17568 21107 17574
rect 21213 17568 21216 17574
rect 21104 17554 21216 17568
rect 21104 17548 21107 17554
rect 21213 17548 21216 17554
rect 21242 17568 21245 17574
rect 22455 17568 22458 17574
rect 21242 17554 22458 17568
rect 21242 17548 21245 17554
rect 22455 17548 22458 17554
rect 22484 17548 22487 17574
rect 25523 17568 25537 17622
rect 25768 17620 25774 17637
rect 25791 17636 25797 17637
rect 27239 17636 27242 17642
rect 25791 17622 27242 17636
rect 25791 17620 25797 17622
rect 25768 17617 25797 17620
rect 27239 17616 27242 17622
rect 27268 17616 27271 17642
rect 26135 17582 26138 17608
rect 26164 17602 26167 17608
rect 26319 17602 26322 17608
rect 26164 17588 26322 17602
rect 26164 17582 26167 17588
rect 26319 17582 26322 17588
rect 26348 17602 26351 17608
rect 26917 17602 26920 17608
rect 26348 17588 26920 17602
rect 26348 17582 26351 17588
rect 26917 17582 26920 17588
rect 26946 17582 26949 17608
rect 25523 17554 28044 17568
rect 19954 17520 20707 17534
rect 22617 17535 22646 17538
rect 19954 17514 19957 17520
rect 22617 17518 22623 17535
rect 22640 17534 22646 17535
rect 22777 17534 22780 17540
rect 22640 17520 22780 17534
rect 22640 17518 22646 17520
rect 22617 17515 22646 17518
rect 22777 17514 22780 17520
rect 22806 17534 22809 17540
rect 23099 17534 23102 17540
rect 22806 17520 23102 17534
rect 22806 17514 22809 17520
rect 23099 17514 23102 17520
rect 23128 17514 23131 17540
rect 24157 17514 24160 17540
rect 24186 17534 24189 17540
rect 24433 17534 24436 17540
rect 24186 17520 24436 17534
rect 24186 17514 24189 17520
rect 24433 17514 24436 17520
rect 24462 17534 24465 17540
rect 24480 17535 24509 17538
rect 24480 17534 24486 17535
rect 24462 17520 24486 17534
rect 24462 17514 24465 17520
rect 24480 17518 24486 17520
rect 24503 17518 24509 17535
rect 24480 17515 24509 17518
rect 24617 17514 24620 17540
rect 24646 17538 24649 17540
rect 24646 17535 24670 17538
rect 24646 17518 24647 17535
rect 24664 17534 24670 17535
rect 25629 17534 25632 17540
rect 24664 17520 25632 17534
rect 24664 17518 24670 17520
rect 24646 17515 24670 17518
rect 24646 17514 24649 17515
rect 25629 17514 25632 17520
rect 25658 17514 25661 17540
rect 25767 17514 25770 17540
rect 25796 17514 25799 17540
rect 25868 17538 25882 17554
rect 26089 17538 26092 17540
rect 25845 17535 25882 17538
rect 25845 17518 25851 17535
rect 25868 17520 25882 17535
rect 25926 17535 25955 17538
rect 25868 17518 25874 17520
rect 25845 17515 25874 17518
rect 25926 17518 25932 17535
rect 25949 17518 25955 17535
rect 26029 17535 26058 17538
rect 25926 17515 25955 17518
rect 25974 17525 26003 17528
rect 21627 17500 21630 17506
rect 19313 17486 21630 17500
rect 19097 17466 19100 17472
rect 18784 17452 19100 17466
rect 19097 17446 19100 17452
rect 19126 17466 19129 17472
rect 19313 17466 19327 17486
rect 21627 17480 21630 17486
rect 21656 17500 21659 17506
rect 22041 17500 22044 17506
rect 21656 17486 22044 17500
rect 21656 17480 21659 17486
rect 22041 17480 22044 17486
rect 22070 17480 22073 17506
rect 22685 17504 22688 17506
rect 22667 17501 22688 17504
rect 22667 17484 22673 17501
rect 22667 17481 22688 17484
rect 22685 17480 22688 17481
rect 22714 17480 22717 17506
rect 24525 17480 24528 17506
rect 24554 17500 24557 17506
rect 24687 17501 24716 17504
rect 24687 17500 24693 17501
rect 24554 17486 24693 17500
rect 24554 17480 24557 17486
rect 24687 17484 24693 17486
rect 24710 17484 24716 17501
rect 24687 17481 24716 17484
rect 25515 17501 25544 17504
rect 25515 17484 25521 17501
rect 25538 17500 25544 17501
rect 25927 17500 25941 17515
rect 25974 17508 25980 17525
rect 25997 17508 26003 17525
rect 26029 17518 26035 17535
rect 26052 17534 26058 17535
rect 26080 17535 26092 17538
rect 26052 17518 26066 17534
rect 26029 17515 26066 17518
rect 26080 17518 26086 17535
rect 26080 17515 26092 17518
rect 25974 17505 26003 17508
rect 25538 17486 25941 17500
rect 25538 17484 25544 17486
rect 25515 17481 25544 17484
rect 19126 17452 19327 17466
rect 19126 17446 19129 17452
rect 25859 17446 25862 17472
rect 25888 17466 25891 17472
rect 25975 17466 25989 17505
rect 26052 17500 26066 17515
rect 26089 17514 26092 17515
rect 26118 17514 26121 17540
rect 26181 17514 26184 17540
rect 26210 17534 26213 17540
rect 26733 17534 26736 17540
rect 26210 17520 26736 17534
rect 26210 17514 26213 17520
rect 26733 17514 26736 17520
rect 26762 17534 26765 17540
rect 27975 17534 27978 17540
rect 26762 17520 27978 17534
rect 26762 17514 26765 17520
rect 27975 17514 27978 17520
rect 28004 17514 28007 17540
rect 28030 17534 28044 17554
rect 29585 17534 29588 17540
rect 28030 17520 29588 17534
rect 29585 17514 29588 17520
rect 29614 17514 29617 17540
rect 26365 17500 26368 17506
rect 26052 17486 26368 17500
rect 26365 17480 26368 17486
rect 26394 17480 26397 17506
rect 28021 17480 28024 17506
rect 28050 17500 28053 17506
rect 28205 17504 28208 17506
rect 28136 17501 28165 17504
rect 28136 17500 28142 17501
rect 28050 17486 28142 17500
rect 28050 17480 28053 17486
rect 28136 17484 28142 17486
rect 28159 17484 28165 17501
rect 28136 17481 28165 17484
rect 28187 17501 28208 17504
rect 28187 17484 28193 17501
rect 28187 17481 28208 17484
rect 28205 17480 28208 17481
rect 28234 17480 28237 17506
rect 25888 17452 25989 17466
rect 29011 17467 29040 17470
rect 25888 17446 25891 17452
rect 29011 17450 29017 17467
rect 29034 17466 29040 17467
rect 29493 17466 29496 17472
rect 29034 17452 29496 17466
rect 29034 17450 29040 17452
rect 29011 17447 29040 17450
rect 29493 17446 29496 17452
rect 29522 17446 29525 17472
rect 3036 17384 29992 17432
rect 4631 17365 4660 17368
rect 4631 17348 4637 17365
rect 4654 17364 4660 17365
rect 4791 17364 4794 17370
rect 4654 17350 4794 17364
rect 4654 17348 4660 17350
rect 4631 17345 4660 17348
rect 4791 17344 4794 17350
rect 4820 17344 4823 17370
rect 18753 17365 18782 17368
rect 18753 17348 18759 17365
rect 18776 17364 18782 17365
rect 18913 17364 18916 17370
rect 18776 17350 18916 17364
rect 18776 17348 18782 17350
rect 18753 17345 18782 17348
rect 18913 17344 18916 17350
rect 18942 17344 18945 17370
rect 26365 17344 26368 17370
rect 26394 17368 26397 17370
rect 26394 17365 26418 17368
rect 26394 17348 26395 17365
rect 26412 17348 26418 17365
rect 27331 17364 27334 17370
rect 26394 17345 26418 17348
rect 26394 17344 26397 17345
rect 27323 17344 27334 17364
rect 27360 17344 27363 17370
rect 3825 17334 3828 17336
rect 3807 17331 3828 17334
rect 3006 17316 3066 17330
rect 3052 17296 3066 17316
rect 3807 17314 3813 17331
rect 3807 17311 3828 17314
rect 3825 17310 3828 17311
rect 3854 17310 3857 17336
rect 7459 17334 7462 17336
rect 7441 17331 7462 17334
rect 7441 17314 7447 17331
rect 7441 17311 7462 17314
rect 7459 17310 7462 17311
rect 7488 17310 7491 17336
rect 12611 17310 12614 17336
rect 12640 17330 12643 17336
rect 12841 17334 12844 17336
rect 12823 17331 12844 17334
rect 12823 17330 12829 17331
rect 12640 17316 12829 17330
rect 12640 17310 12643 17316
rect 12823 17314 12829 17316
rect 12823 17311 12844 17314
rect 12841 17310 12844 17311
rect 12870 17310 12873 17336
rect 14451 17310 14454 17336
rect 14480 17330 14483 17336
rect 14881 17331 14910 17334
rect 14881 17330 14887 17331
rect 14480 17316 14887 17330
rect 14480 17310 14483 17316
rect 14881 17314 14887 17316
rect 14904 17314 14910 17331
rect 14881 17311 14910 17314
rect 17929 17331 17958 17334
rect 17929 17314 17935 17331
rect 17952 17330 17958 17331
rect 17993 17330 17996 17336
rect 17952 17316 17996 17330
rect 17952 17314 17958 17316
rect 17929 17311 17958 17314
rect 17993 17310 17996 17316
rect 18022 17310 18025 17336
rect 20459 17331 20488 17334
rect 20459 17314 20465 17331
rect 20482 17330 20488 17331
rect 23173 17331 23202 17334
rect 20482 17316 20592 17330
rect 20482 17314 20488 17316
rect 20459 17311 20488 17314
rect 3757 17297 3786 17300
rect 3757 17296 3763 17297
rect 3052 17282 3763 17296
rect 3757 17280 3763 17282
rect 3780 17296 3786 17297
rect 5757 17296 5760 17302
rect 3780 17282 5760 17296
rect 3780 17280 3786 17282
rect 3757 17277 3786 17280
rect 5757 17276 5760 17282
rect 5786 17276 5789 17302
rect 6953 17276 6956 17302
rect 6982 17296 6985 17302
rect 7229 17296 7232 17302
rect 6982 17282 7232 17296
rect 6982 17276 6985 17282
rect 7229 17276 7232 17282
rect 7258 17276 7261 17302
rect 7391 17297 7420 17300
rect 7391 17280 7397 17297
rect 7414 17296 7420 17297
rect 7551 17296 7554 17302
rect 7414 17282 7554 17296
rect 7414 17280 7420 17282
rect 7391 17277 7420 17280
rect 7551 17276 7554 17282
rect 7580 17296 7583 17302
rect 7873 17296 7876 17302
rect 7580 17282 7876 17296
rect 7580 17276 7583 17282
rect 7873 17276 7876 17282
rect 7902 17276 7905 17302
rect 12657 17276 12660 17302
rect 12686 17276 12689 17302
rect 12773 17297 12802 17300
rect 12773 17280 12779 17297
rect 12796 17296 12802 17297
rect 12933 17296 12936 17302
rect 12796 17282 12936 17296
rect 12796 17280 12802 17282
rect 12773 17277 12802 17280
rect 12933 17276 12936 17282
rect 12962 17276 12965 17302
rect 13945 17276 13948 17302
rect 13974 17296 13977 17302
rect 14837 17297 14866 17300
rect 14837 17296 14843 17297
rect 13974 17282 14843 17296
rect 13974 17276 13977 17282
rect 14837 17280 14843 17282
rect 14860 17280 14866 17297
rect 14837 17277 14866 17280
rect 17717 17276 17720 17302
rect 17746 17276 17749 17302
rect 17855 17276 17858 17302
rect 17884 17300 17887 17302
rect 17884 17297 17902 17300
rect 17896 17280 17902 17297
rect 18002 17296 18016 17310
rect 19649 17296 19652 17302
rect 18002 17282 19652 17296
rect 17884 17277 17902 17280
rect 17884 17276 17887 17277
rect 19649 17276 19652 17282
rect 19678 17276 19681 17302
rect 20155 17276 20158 17302
rect 20184 17296 20187 17302
rect 20403 17297 20432 17300
rect 20403 17296 20409 17297
rect 20184 17282 20409 17296
rect 20184 17276 20187 17282
rect 20403 17280 20409 17282
rect 20426 17280 20432 17297
rect 20578 17296 20592 17316
rect 23173 17314 23179 17331
rect 23196 17330 23202 17331
rect 23237 17330 23240 17336
rect 23196 17316 23240 17330
rect 23196 17314 23202 17316
rect 23173 17311 23202 17314
rect 23237 17310 23240 17316
rect 23266 17310 23269 17336
rect 25583 17334 25586 17336
rect 25565 17331 25586 17334
rect 25565 17314 25571 17331
rect 25565 17311 25586 17314
rect 25583 17310 25586 17311
rect 25612 17310 25615 17336
rect 27055 17310 27058 17336
rect 27084 17330 27087 17336
rect 27084 17316 27170 17330
rect 27084 17310 27087 17316
rect 20799 17296 20802 17302
rect 20578 17282 20802 17296
rect 20403 17277 20432 17280
rect 20799 17276 20802 17282
rect 20828 17276 20831 17302
rect 23099 17276 23102 17302
rect 23128 17300 23131 17302
rect 23128 17297 23146 17300
rect 23140 17280 23146 17297
rect 23128 17277 23146 17280
rect 25515 17297 25544 17300
rect 25515 17280 25521 17297
rect 25538 17296 25544 17297
rect 25629 17296 25632 17302
rect 25538 17282 25632 17296
rect 25538 17280 25544 17282
rect 25515 17277 25544 17280
rect 23128 17276 23131 17277
rect 25629 17276 25632 17282
rect 25658 17276 25661 17302
rect 27101 17276 27104 17302
rect 27130 17276 27133 17302
rect 27156 17300 27170 17316
rect 27323 17311 27337 17344
rect 28435 17334 28438 17336
rect 28417 17331 28438 17334
rect 28417 17314 28423 17331
rect 28417 17311 28438 17314
rect 27315 17308 27344 17311
rect 28435 17310 28438 17311
rect 28464 17310 28467 17336
rect 29493 17310 29496 17336
rect 29522 17310 29525 17336
rect 27156 17297 27188 17300
rect 27156 17282 27165 17297
rect 27159 17280 27165 17282
rect 27182 17280 27188 17297
rect 27159 17277 27188 17280
rect 27239 17276 27242 17302
rect 27268 17300 27271 17302
rect 27268 17297 27289 17300
rect 27283 17280 27289 17297
rect 27315 17291 27321 17308
rect 27338 17291 27344 17308
rect 27423 17300 27426 17302
rect 27315 17288 27344 17291
rect 27363 17297 27392 17300
rect 27268 17277 27289 17280
rect 27363 17280 27369 17297
rect 27386 17280 27392 17297
rect 27363 17277 27392 17280
rect 27414 17297 27426 17300
rect 27414 17280 27420 17297
rect 27414 17277 27426 17280
rect 27268 17276 27271 17277
rect 3135 17242 3138 17268
rect 3164 17262 3167 17268
rect 3596 17263 3625 17266
rect 3596 17262 3602 17263
rect 3164 17248 3602 17262
rect 3164 17242 3167 17248
rect 3596 17246 3602 17248
rect 3619 17246 3625 17263
rect 3596 17243 3625 17246
rect 12612 17263 12641 17266
rect 12612 17246 12618 17263
rect 12635 17262 12641 17263
rect 12666 17262 12680 17276
rect 12635 17248 12680 17262
rect 12635 17246 12641 17248
rect 12612 17243 12641 17246
rect 8425 17208 8428 17234
rect 8454 17228 8457 17234
rect 8655 17228 8658 17234
rect 8454 17214 8658 17228
rect 8454 17208 8457 17214
rect 8655 17208 8658 17214
rect 8684 17228 8687 17234
rect 10035 17228 10038 17234
rect 8684 17214 10038 17228
rect 8684 17208 8687 17214
rect 10035 17208 10038 17214
rect 10064 17228 10067 17234
rect 10173 17228 10176 17234
rect 10064 17214 10176 17228
rect 10064 17208 10067 17214
rect 10173 17208 10176 17214
rect 10202 17228 10205 17234
rect 10587 17228 10590 17234
rect 10202 17214 10590 17228
rect 10202 17208 10205 17214
rect 10587 17208 10590 17214
rect 10616 17228 10619 17234
rect 10909 17228 10912 17234
rect 10616 17214 10912 17228
rect 10616 17208 10619 17214
rect 10909 17208 10912 17214
rect 10938 17228 10941 17234
rect 12620 17228 12634 17243
rect 14497 17242 14500 17268
rect 14526 17262 14529 17268
rect 14682 17263 14711 17266
rect 14682 17262 14688 17263
rect 14526 17248 14688 17262
rect 14526 17242 14529 17248
rect 14682 17246 14688 17248
rect 14705 17246 14711 17263
rect 14682 17243 14711 17246
rect 17027 17242 17030 17268
rect 17056 17262 17059 17268
rect 17671 17262 17674 17268
rect 17056 17248 17674 17262
rect 17056 17242 17059 17248
rect 17671 17242 17674 17248
rect 17700 17242 17703 17268
rect 20248 17263 20277 17266
rect 20248 17246 20254 17263
rect 20271 17246 20277 17263
rect 20248 17243 20277 17246
rect 22962 17263 22991 17266
rect 22962 17246 22968 17263
rect 22985 17246 22991 17263
rect 22962 17243 22991 17246
rect 10938 17214 12634 17228
rect 10938 17208 10941 17214
rect 8287 17198 8290 17200
rect 8265 17195 8290 17198
rect 8265 17178 8271 17195
rect 8288 17178 8290 17195
rect 8265 17175 8290 17178
rect 8287 17174 8290 17175
rect 8316 17174 8319 17200
rect 9621 17174 9624 17200
rect 9650 17194 9653 17200
rect 11645 17194 11648 17200
rect 9650 17180 11648 17194
rect 9650 17174 9653 17180
rect 11645 17174 11648 17180
rect 11674 17174 11677 17200
rect 13647 17195 13676 17198
rect 13647 17178 13653 17195
rect 13670 17194 13676 17195
rect 14313 17194 14316 17200
rect 13670 17180 14316 17194
rect 13670 17178 13676 17180
rect 13647 17175 13676 17178
rect 14313 17174 14316 17180
rect 14342 17174 14345 17200
rect 15233 17174 15236 17200
rect 15262 17194 15265 17200
rect 15717 17195 15746 17198
rect 15717 17194 15723 17195
rect 15262 17180 15723 17194
rect 15262 17174 15265 17180
rect 15717 17178 15723 17180
rect 15740 17178 15746 17195
rect 20256 17194 20270 17243
rect 20569 17194 20572 17200
rect 20256 17180 20572 17194
rect 15717 17175 15746 17178
rect 20569 17174 20572 17180
rect 20598 17174 20601 17200
rect 21283 17195 21312 17198
rect 21283 17178 21289 17195
rect 21306 17194 21312 17195
rect 21443 17194 21446 17200
rect 21306 17180 21446 17194
rect 21306 17178 21312 17180
rect 21283 17175 21312 17178
rect 21443 17174 21446 17180
rect 21472 17174 21475 17200
rect 22970 17194 22984 17243
rect 24709 17242 24712 17268
rect 24738 17262 24741 17268
rect 25354 17263 25383 17266
rect 25354 17262 25360 17263
rect 24738 17248 25360 17262
rect 24738 17242 24741 17248
rect 25354 17246 25360 17248
rect 25377 17246 25383 17263
rect 27371 17262 27385 17277
rect 27423 17276 27426 17277
rect 27452 17276 27455 17302
rect 28021 17296 28024 17302
rect 27800 17282 28024 17296
rect 27745 17262 27748 17268
rect 27371 17248 27748 17262
rect 25354 17243 25383 17246
rect 23997 17229 24026 17232
rect 23997 17212 24003 17229
rect 24020 17228 24026 17229
rect 24295 17228 24298 17234
rect 24020 17214 24298 17228
rect 24020 17212 24026 17214
rect 23997 17209 24026 17212
rect 24295 17208 24298 17214
rect 24324 17208 24327 17234
rect 23145 17194 23148 17200
rect 22970 17180 23148 17194
rect 23145 17174 23148 17180
rect 23174 17174 23177 17200
rect 25362 17194 25376 17243
rect 27745 17242 27748 17248
rect 27774 17242 27777 17268
rect 26779 17208 26782 17234
rect 26808 17228 26811 17234
rect 27800 17228 27814 17282
rect 28021 17276 28024 17282
rect 28050 17296 28053 17302
rect 28343 17296 28346 17302
rect 28372 17300 28375 17302
rect 28372 17297 28390 17300
rect 28050 17282 28346 17296
rect 28050 17276 28053 17282
rect 28343 17276 28346 17282
rect 28384 17280 28390 17297
rect 28372 17277 28390 17280
rect 28372 17276 28375 17277
rect 29401 17276 29404 17302
rect 29430 17296 29433 17302
rect 29586 17297 29615 17300
rect 29586 17296 29592 17297
rect 29430 17282 29592 17296
rect 29430 17276 29433 17282
rect 29586 17280 29592 17282
rect 29609 17280 29615 17297
rect 29586 17277 29615 17280
rect 29632 17297 29661 17300
rect 29632 17280 29638 17297
rect 29655 17280 29661 17297
rect 29632 17277 29661 17280
rect 29696 17297 29725 17300
rect 29696 17280 29702 17297
rect 29719 17296 29725 17297
rect 29769 17296 29772 17302
rect 29719 17282 29772 17296
rect 29719 17280 29725 17282
rect 29696 17277 29725 17280
rect 27975 17242 27978 17268
rect 28004 17262 28007 17268
rect 28206 17263 28235 17266
rect 28206 17262 28212 17263
rect 28004 17248 28212 17262
rect 28004 17242 28007 17248
rect 28206 17246 28212 17248
rect 28229 17246 28235 17263
rect 28206 17243 28235 17246
rect 29241 17263 29270 17266
rect 29241 17246 29247 17263
rect 29264 17262 29270 17263
rect 29640 17262 29654 17277
rect 29769 17276 29772 17282
rect 29798 17276 29801 17302
rect 29264 17248 29654 17262
rect 29264 17246 29270 17248
rect 29241 17243 29270 17246
rect 26808 17214 27814 17228
rect 26808 17208 26811 17214
rect 26733 17194 26736 17200
rect 25362 17180 26736 17194
rect 26733 17174 26736 17180
rect 26762 17174 26765 17200
rect 27102 17195 27131 17198
rect 27102 17178 27108 17195
rect 27125 17194 27131 17195
rect 28619 17194 28622 17200
rect 27125 17180 28622 17194
rect 27125 17178 27131 17180
rect 27102 17175 27131 17178
rect 28619 17174 28622 17180
rect 28648 17174 28651 17200
rect 29493 17174 29496 17200
rect 29522 17174 29525 17200
rect 3036 17112 29992 17160
rect 5665 17092 5668 17098
rect 5490 17078 5668 17092
rect 5490 17028 5504 17078
rect 5665 17072 5668 17078
rect 5694 17072 5697 17098
rect 6517 17093 6546 17096
rect 6517 17076 6523 17093
rect 6540 17092 6546 17093
rect 6677 17092 6680 17098
rect 6540 17078 6680 17092
rect 6540 17076 6546 17078
rect 6517 17073 6546 17076
rect 6677 17072 6680 17078
rect 6706 17072 6709 17098
rect 11967 17092 11970 17098
rect 9538 17078 11970 17092
rect 5482 17025 5511 17028
rect 5482 17008 5488 17025
rect 5505 17008 5511 17025
rect 5482 17005 5511 17008
rect 8655 17004 8658 17030
rect 8684 17004 8687 17030
rect 5643 16991 5672 16994
rect 5643 16974 5649 16991
rect 5666 16990 5672 16991
rect 5757 16990 5760 16996
rect 5666 16976 5760 16990
rect 5666 16974 5672 16976
rect 5643 16971 5672 16974
rect 5757 16970 5760 16976
rect 5786 16970 5789 16996
rect 6079 16990 6082 16996
rect 5812 16976 6082 16990
rect 5693 16957 5722 16960
rect 5693 16940 5699 16957
rect 5716 16956 5722 16957
rect 5812 16956 5826 16976
rect 6079 16970 6082 16976
rect 6108 16990 6111 16996
rect 7045 16990 7048 16996
rect 6108 16976 7048 16990
rect 6108 16970 6111 16976
rect 7045 16970 7048 16976
rect 7074 16970 7077 16996
rect 8817 16991 8846 16994
rect 8817 16974 8823 16991
rect 8840 16990 8846 16991
rect 8977 16990 8980 16996
rect 8840 16976 8980 16990
rect 8840 16974 8846 16976
rect 8817 16971 8846 16974
rect 8977 16970 8980 16976
rect 9006 16990 9009 16996
rect 9538 16990 9552 17078
rect 11967 17072 11970 17078
rect 11996 17072 11999 17098
rect 24433 17072 24436 17098
rect 24462 17092 24465 17098
rect 24709 17092 24712 17098
rect 24462 17078 24712 17092
rect 24462 17072 24465 17078
rect 10909 17004 10912 17030
rect 10938 17024 10941 17030
rect 10956 17025 10985 17028
rect 10956 17024 10962 17025
rect 10938 17010 10962 17024
rect 10938 17004 10941 17010
rect 10956 17008 10962 17010
rect 10979 17008 10985 17025
rect 10956 17005 10985 17008
rect 11991 17025 12020 17028
rect 11991 17008 11997 17025
rect 12014 17024 12020 17025
rect 12014 17010 12358 17024
rect 12014 17008 12020 17010
rect 11991 17005 12020 17008
rect 9006 16976 9552 16990
rect 9006 16970 9009 16976
rect 12243 16970 12246 16996
rect 12272 16970 12275 16996
rect 12344 16994 12358 17010
rect 12749 17004 12752 17030
rect 12778 17024 12781 17030
rect 12934 17025 12963 17028
rect 12934 17024 12940 17025
rect 12778 17010 12940 17024
rect 12778 17004 12781 17010
rect 12934 17008 12940 17010
rect 12957 17008 12963 17025
rect 12934 17005 12963 17008
rect 14774 17025 14803 17028
rect 14774 17008 14780 17025
rect 14797 17024 14803 17025
rect 15003 17024 15006 17030
rect 14797 17010 15006 17024
rect 14797 17008 14803 17010
rect 14774 17005 14803 17008
rect 15003 17004 15006 17010
rect 15032 17004 15035 17030
rect 21213 17024 21216 17030
rect 15150 17010 15854 17024
rect 15150 16996 15164 17010
rect 12336 16991 12365 16994
rect 12336 16974 12342 16991
rect 12359 16974 12365 16991
rect 12336 16971 12365 16974
rect 14727 16970 14730 16996
rect 14756 16970 14759 16996
rect 14838 16991 14867 16994
rect 14838 16974 14844 16991
rect 14861 16990 14867 16991
rect 14861 16976 15118 16990
rect 14861 16974 14867 16976
rect 14838 16971 14867 16974
rect 5716 16942 5826 16956
rect 5716 16940 5722 16942
rect 5693 16937 5722 16940
rect 7137 16936 7140 16962
rect 7166 16956 7169 16962
rect 7459 16956 7462 16962
rect 7166 16942 7462 16956
rect 7166 16936 7169 16942
rect 7459 16936 7462 16942
rect 7488 16956 7491 16962
rect 8863 16957 8892 16960
rect 8863 16956 8869 16957
rect 7488 16942 8869 16956
rect 7488 16936 7491 16942
rect 8863 16940 8869 16942
rect 8886 16956 8892 16957
rect 8931 16956 8934 16962
rect 8886 16942 8934 16956
rect 8886 16940 8892 16942
rect 8863 16937 8892 16940
rect 8931 16936 8934 16942
rect 8960 16936 8963 16962
rect 10127 16936 10130 16962
rect 10156 16956 10159 16962
rect 10633 16956 10636 16962
rect 10156 16942 10636 16956
rect 10156 16936 10159 16942
rect 10633 16936 10636 16942
rect 10662 16956 10665 16962
rect 11185 16960 11188 16962
rect 11116 16957 11145 16960
rect 11116 16956 11122 16957
rect 10662 16942 11122 16956
rect 10662 16936 10665 16942
rect 11116 16940 11122 16942
rect 11139 16940 11145 16957
rect 11116 16937 11145 16940
rect 11167 16957 11188 16960
rect 11167 16940 11173 16957
rect 11167 16937 11188 16940
rect 11185 16936 11188 16937
rect 11214 16936 11217 16962
rect 12933 16936 12936 16962
rect 12962 16956 12965 16962
rect 13163 16960 13166 16962
rect 13094 16957 13123 16960
rect 13094 16956 13100 16957
rect 12962 16942 13100 16956
rect 12962 16936 12965 16942
rect 13094 16940 13100 16942
rect 13117 16940 13123 16957
rect 13094 16937 13123 16940
rect 13145 16957 13166 16960
rect 13145 16940 13151 16957
rect 13145 16937 13166 16940
rect 13163 16936 13166 16937
rect 13192 16936 13195 16962
rect 14037 16936 14040 16962
rect 14066 16956 14069 16962
rect 14636 16957 14665 16960
rect 14636 16956 14642 16957
rect 14066 16942 14642 16956
rect 14066 16936 14069 16942
rect 14636 16940 14642 16942
rect 14659 16940 14665 16957
rect 14636 16937 14665 16940
rect 14773 16936 14776 16962
rect 14802 16936 14805 16962
rect 15104 16956 15118 16976
rect 15141 16970 15144 16996
rect 15170 16970 15173 16996
rect 15233 16970 15236 16996
rect 15262 16970 15265 16996
rect 15463 16970 15466 16996
rect 15492 16990 15495 16996
rect 15786 16991 15815 16994
rect 15786 16990 15792 16991
rect 15492 16976 15792 16990
rect 15492 16970 15495 16976
rect 15786 16974 15792 16976
rect 15809 16974 15815 16991
rect 15840 16990 15854 17010
rect 20693 17010 21216 17024
rect 17074 16991 17103 16994
rect 16024 16990 16084 16991
rect 17074 16990 17080 16991
rect 15840 16977 17080 16990
rect 15840 16976 16038 16977
rect 16070 16976 17080 16977
rect 15786 16971 15815 16974
rect 17074 16974 17080 16976
rect 17097 16990 17103 16991
rect 17119 16990 17122 16996
rect 17097 16976 17122 16990
rect 17097 16974 17103 16976
rect 17074 16971 17103 16974
rect 17119 16970 17122 16976
rect 17148 16970 17151 16996
rect 17165 16970 17168 16996
rect 17194 16970 17197 16996
rect 20569 16970 20572 16996
rect 20598 16990 20601 16996
rect 20693 16990 20707 17010
rect 21213 17004 21216 17010
rect 21242 17004 21245 17030
rect 24534 17028 24548 17078
rect 24709 17072 24712 17078
rect 24738 17072 24741 17098
rect 25561 17093 25590 17096
rect 25561 17076 25567 17093
rect 25584 17092 25590 17093
rect 25767 17092 25770 17098
rect 25584 17078 25770 17092
rect 25584 17076 25590 17078
rect 25561 17073 25590 17076
rect 25767 17072 25770 17078
rect 25796 17072 25799 17098
rect 26135 17072 26138 17098
rect 26164 17092 26167 17098
rect 26963 17092 26966 17098
rect 26164 17078 26966 17092
rect 26164 17072 26167 17078
rect 26963 17072 26966 17078
rect 26992 17072 26995 17098
rect 27745 17072 27748 17098
rect 27774 17096 27777 17098
rect 27774 17093 27798 17096
rect 27774 17076 27775 17093
rect 27792 17076 27798 17093
rect 27774 17073 27798 17076
rect 27774 17072 27777 17073
rect 27975 17072 27978 17098
rect 28004 17092 28007 17098
rect 28389 17092 28392 17098
rect 28004 17078 28392 17092
rect 28004 17072 28007 17078
rect 28389 17072 28392 17078
rect 28418 17072 28421 17098
rect 24526 17025 24555 17028
rect 24526 17008 24532 17025
rect 24549 17008 24555 17025
rect 24526 17005 24555 17008
rect 25523 17010 26802 17024
rect 20598 16976 20707 16990
rect 21375 16991 21404 16994
rect 20598 16970 20601 16976
rect 21375 16974 21381 16991
rect 21398 16990 21404 16991
rect 21489 16990 21492 16996
rect 21398 16976 21492 16990
rect 21398 16974 21404 16976
rect 21375 16971 21404 16974
rect 21489 16970 21492 16976
rect 21518 16970 21521 16996
rect 21535 16970 21538 16996
rect 21564 16970 21567 16996
rect 24571 16970 24574 16996
rect 24600 16990 24603 16996
rect 24681 16991 24710 16994
rect 24681 16990 24687 16991
rect 24600 16976 24687 16990
rect 24600 16970 24603 16976
rect 24681 16974 24687 16976
rect 24704 16974 24710 16991
rect 25523 16990 25537 17010
rect 24681 16971 24710 16974
rect 24856 16976 25537 16990
rect 15647 16956 15650 16962
rect 15104 16942 15650 16956
rect 15647 16936 15650 16942
rect 15676 16936 15679 16962
rect 15831 16936 15834 16962
rect 15860 16956 15863 16962
rect 16015 16960 16018 16962
rect 15946 16957 15975 16960
rect 15946 16956 15952 16957
rect 15860 16942 15952 16956
rect 15860 16936 15863 16942
rect 15946 16940 15952 16942
rect 15969 16940 15975 16957
rect 15946 16937 15975 16940
rect 15997 16957 16018 16960
rect 15997 16940 16003 16957
rect 15997 16937 16018 16940
rect 16015 16936 16018 16937
rect 16044 16936 16047 16962
rect 21425 16957 21454 16960
rect 21425 16940 21431 16957
rect 21448 16956 21454 16957
rect 21544 16956 21558 16970
rect 21448 16942 21558 16956
rect 21448 16940 21454 16942
rect 21425 16937 21454 16940
rect 22685 16936 22688 16962
rect 22714 16956 22717 16962
rect 24725 16957 24754 16960
rect 24725 16956 24731 16957
rect 22714 16942 24731 16956
rect 22714 16936 22717 16942
rect 24725 16940 24731 16942
rect 24748 16956 24754 16957
rect 24856 16956 24870 16976
rect 26733 16970 26736 16996
rect 26762 16970 26765 16996
rect 26788 16990 26802 17010
rect 28619 17004 28622 17030
rect 28648 17004 28651 17030
rect 28297 16990 28300 16996
rect 26788 16976 28300 16990
rect 28297 16970 28300 16976
rect 28326 16970 28329 16996
rect 28712 16991 28741 16994
rect 28712 16974 28718 16991
rect 28735 16990 28741 16991
rect 29493 16990 29496 16996
rect 28735 16976 29496 16990
rect 28735 16974 28741 16976
rect 28712 16971 28741 16974
rect 29493 16970 29496 16976
rect 29522 16970 29525 16996
rect 24748 16942 24870 16956
rect 24748 16940 24754 16942
rect 24725 16937 24754 16940
rect 26411 16936 26414 16962
rect 26440 16956 26443 16962
rect 26779 16956 26782 16962
rect 26440 16942 26782 16956
rect 26440 16936 26443 16942
rect 26779 16936 26782 16942
rect 26808 16956 26811 16962
rect 26963 16960 26966 16962
rect 26895 16957 26924 16960
rect 26895 16956 26901 16957
rect 26808 16942 26901 16956
rect 26808 16936 26811 16942
rect 26895 16940 26901 16942
rect 26918 16940 26924 16957
rect 26895 16937 26924 16940
rect 26945 16957 26966 16960
rect 26945 16940 26951 16957
rect 26945 16937 26966 16940
rect 26963 16936 26966 16937
rect 26992 16936 26995 16962
rect 28804 16957 28833 16960
rect 28804 16940 28810 16957
rect 28827 16940 28833 16957
rect 28804 16937 28833 16940
rect 9529 16902 9532 16928
rect 9558 16922 9561 16928
rect 9691 16923 9720 16926
rect 9691 16922 9697 16923
rect 9558 16908 9697 16922
rect 9558 16902 9561 16908
rect 9691 16906 9697 16908
rect 9714 16906 9720 16923
rect 9691 16903 9720 16906
rect 12105 16902 12108 16928
rect 12134 16922 12137 16928
rect 12290 16923 12319 16926
rect 12290 16922 12296 16923
rect 12134 16908 12296 16922
rect 12134 16902 12137 16908
rect 12290 16906 12296 16908
rect 12313 16906 12319 16923
rect 12290 16903 12319 16906
rect 13969 16923 13998 16926
rect 13969 16906 13975 16923
rect 13992 16922 13998 16923
rect 14267 16922 14270 16928
rect 13992 16908 14270 16922
rect 13992 16906 13998 16908
rect 13969 16903 13998 16906
rect 14267 16902 14270 16908
rect 14296 16902 14299 16928
rect 14865 16902 14868 16928
rect 14894 16922 14897 16928
rect 15188 16923 15217 16926
rect 15188 16922 15194 16923
rect 14894 16908 15194 16922
rect 14894 16902 14897 16908
rect 15188 16906 15194 16908
rect 15211 16906 15217 16923
rect 15188 16903 15217 16906
rect 16821 16923 16850 16926
rect 16821 16906 16827 16923
rect 16844 16922 16850 16923
rect 17073 16922 17076 16928
rect 16844 16908 17076 16922
rect 16844 16906 16850 16908
rect 16821 16903 16850 16906
rect 17073 16902 17076 16908
rect 17102 16902 17105 16928
rect 17166 16923 17195 16926
rect 17166 16906 17172 16923
rect 17189 16922 17195 16923
rect 17303 16922 17306 16928
rect 17189 16908 17306 16922
rect 17189 16906 17195 16908
rect 17166 16903 17195 16906
rect 17303 16902 17306 16908
rect 17332 16902 17335 16928
rect 21673 16902 21676 16928
rect 21702 16922 21705 16928
rect 22249 16923 22278 16926
rect 22249 16922 22255 16923
rect 21702 16908 22255 16922
rect 21702 16902 21705 16908
rect 22249 16906 22255 16908
rect 22272 16906 22278 16923
rect 22249 16903 22278 16906
rect 28113 16902 28116 16928
rect 28142 16922 28145 16928
rect 28758 16923 28787 16926
rect 28758 16922 28764 16923
rect 28142 16908 28764 16922
rect 28142 16902 28145 16908
rect 28758 16906 28764 16908
rect 28781 16906 28787 16923
rect 28812 16922 28826 16937
rect 28987 16936 28990 16962
rect 29016 16936 29019 16962
rect 29493 16922 29496 16928
rect 28812 16908 29496 16922
rect 28758 16903 28787 16906
rect 29493 16902 29496 16908
rect 29522 16902 29525 16928
rect 3036 16840 29992 16888
rect 13831 16821 13860 16824
rect 13831 16804 13837 16821
rect 13854 16820 13860 16821
rect 14037 16820 14040 16826
rect 13854 16806 14040 16820
rect 13854 16804 13860 16806
rect 13831 16801 13860 16804
rect 14037 16800 14040 16806
rect 14066 16800 14069 16826
rect 14544 16821 14573 16824
rect 14544 16804 14550 16821
rect 14567 16820 14573 16821
rect 14958 16821 14987 16824
rect 14958 16820 14964 16821
rect 14567 16806 14964 16820
rect 14567 16804 14573 16806
rect 14544 16801 14573 16804
rect 14958 16804 14964 16806
rect 14981 16804 14987 16821
rect 14958 16801 14987 16804
rect 15003 16800 15006 16826
rect 15032 16800 15035 16826
rect 15049 16800 15052 16826
rect 15078 16800 15081 16826
rect 18821 16824 18824 16826
rect 18799 16821 18824 16824
rect 18799 16804 18805 16821
rect 18822 16804 18824 16821
rect 18799 16801 18824 16804
rect 18821 16800 18824 16801
rect 18850 16800 18853 16826
rect 21259 16800 21262 16826
rect 21288 16820 21291 16826
rect 21306 16821 21335 16824
rect 21306 16820 21312 16821
rect 21288 16806 21312 16820
rect 21288 16800 21291 16806
rect 21306 16804 21312 16806
rect 21329 16804 21335 16821
rect 21306 16801 21335 16804
rect 22685 16800 22688 16826
rect 22714 16820 22717 16826
rect 23007 16820 23010 16826
rect 22714 16806 23010 16820
rect 22714 16800 22717 16806
rect 23007 16800 23010 16806
rect 23036 16800 23039 16826
rect 27033 16821 27062 16824
rect 27033 16804 27039 16821
rect 27056 16820 27062 16821
rect 27239 16820 27242 16826
rect 27056 16806 27242 16820
rect 27056 16804 27062 16806
rect 27033 16801 27062 16804
rect 27239 16800 27242 16806
rect 27268 16800 27271 16826
rect 7487 16787 7516 16790
rect 7487 16770 7493 16787
rect 7510 16786 7516 16787
rect 7510 16772 7620 16786
rect 7510 16770 7516 16772
rect 7487 16767 7516 16770
rect 7437 16753 7466 16756
rect 7437 16736 7443 16753
rect 7460 16752 7466 16753
rect 7551 16752 7554 16758
rect 7460 16738 7554 16752
rect 7460 16736 7466 16738
rect 7437 16733 7466 16736
rect 7551 16732 7554 16738
rect 7580 16732 7583 16758
rect 7606 16752 7620 16772
rect 8931 16766 8934 16792
rect 8960 16786 8963 16792
rect 10235 16787 10264 16790
rect 10235 16786 10241 16787
rect 8960 16772 10241 16786
rect 8960 16766 8963 16772
rect 10235 16770 10241 16772
rect 10258 16770 10264 16787
rect 10235 16767 10264 16770
rect 11645 16766 11648 16792
rect 11674 16786 11677 16792
rect 12289 16786 12292 16792
rect 11674 16772 12292 16786
rect 11674 16766 11677 16772
rect 12289 16766 12292 16772
rect 12318 16766 12321 16792
rect 12657 16766 12660 16792
rect 12686 16786 12689 16792
rect 13025 16790 13028 16792
rect 13007 16787 13028 16790
rect 13007 16786 13013 16787
rect 12686 16772 13013 16786
rect 12686 16766 12689 16772
rect 13007 16770 13013 16772
rect 13007 16767 13028 16770
rect 13025 16766 13028 16767
rect 13054 16766 13057 16792
rect 14267 16766 14270 16792
rect 14296 16786 14299 16792
rect 14296 16772 14612 16786
rect 14296 16766 14299 16772
rect 8333 16752 8336 16758
rect 7606 16738 8336 16752
rect 8333 16732 8336 16738
rect 8362 16752 8365 16758
rect 8425 16752 8428 16758
rect 8362 16738 8428 16752
rect 8362 16732 8365 16738
rect 8425 16732 8428 16738
rect 8454 16732 8457 16758
rect 9529 16732 9532 16758
rect 9558 16732 9561 16758
rect 9621 16732 9624 16758
rect 9650 16732 9653 16758
rect 9667 16732 9670 16758
rect 9696 16732 9699 16758
rect 9714 16753 9743 16756
rect 9714 16736 9720 16753
rect 9737 16752 9743 16753
rect 9737 16738 9874 16752
rect 9737 16736 9743 16738
rect 9714 16733 9743 16736
rect 7275 16698 7278 16724
rect 7304 16698 7307 16724
rect 8379 16698 8382 16724
rect 8408 16718 8411 16724
rect 9630 16718 9644 16732
rect 8408 16704 9644 16718
rect 8408 16698 8411 16704
rect 9860 16684 9874 16738
rect 10035 16732 10038 16758
rect 10064 16732 10067 16758
rect 10173 16732 10176 16758
rect 10202 16756 10205 16758
rect 10202 16753 10220 16756
rect 10214 16736 10220 16753
rect 10202 16733 10220 16736
rect 11071 16753 11100 16756
rect 11071 16736 11077 16753
rect 11094 16752 11100 16753
rect 11554 16753 11583 16756
rect 11554 16752 11560 16753
rect 11094 16738 11560 16752
rect 11094 16736 11100 16738
rect 11071 16733 11100 16736
rect 11554 16736 11560 16738
rect 11577 16736 11583 16753
rect 11554 16733 11583 16736
rect 10202 16732 10205 16733
rect 11691 16732 11694 16758
rect 11720 16732 11723 16758
rect 11737 16732 11740 16758
rect 11766 16756 11769 16758
rect 11766 16752 11770 16756
rect 12014 16753 12043 16756
rect 11766 16738 11788 16752
rect 11766 16733 11770 16738
rect 12014 16736 12020 16753
rect 12037 16736 12043 16753
rect 12014 16733 12043 16736
rect 11766 16732 11769 16733
rect 11600 16719 11629 16722
rect 11600 16702 11606 16719
rect 11623 16718 11629 16719
rect 12022 16718 12036 16733
rect 12105 16732 12108 16758
rect 12134 16732 12137 16758
rect 12749 16732 12752 16758
rect 12778 16752 12781 16758
rect 12796 16753 12825 16756
rect 12796 16752 12802 16753
rect 12778 16738 12802 16752
rect 12778 16732 12781 16738
rect 12796 16736 12802 16738
rect 12819 16736 12825 16753
rect 12796 16733 12825 16736
rect 12841 16732 12844 16758
rect 12870 16752 12873 16758
rect 12933 16752 12936 16758
rect 12962 16756 12965 16758
rect 12962 16753 12980 16756
rect 12870 16738 12936 16752
rect 12870 16732 12873 16738
rect 12933 16732 12936 16738
rect 12974 16736 12980 16753
rect 12962 16733 12980 16736
rect 12962 16732 12965 16733
rect 14313 16732 14316 16758
rect 14342 16732 14345 16758
rect 14371 16753 14400 16756
rect 14371 16752 14377 16753
rect 14368 16736 14377 16752
rect 14394 16736 14400 16753
rect 14368 16733 14400 16736
rect 11623 16704 12036 16718
rect 11623 16702 11629 16704
rect 11600 16699 11629 16702
rect 13853 16698 13856 16724
rect 13882 16718 13885 16724
rect 14083 16718 14086 16724
rect 13882 16704 14086 16718
rect 13882 16698 13885 16704
rect 14083 16698 14086 16704
rect 14112 16718 14115 16724
rect 14368 16718 14382 16733
rect 14451 16732 14454 16758
rect 14480 16756 14483 16758
rect 14598 16756 14612 16772
rect 14865 16766 14868 16792
rect 14894 16766 14897 16792
rect 15555 16766 15558 16792
rect 15584 16786 15587 16792
rect 15763 16787 15792 16790
rect 15763 16786 15769 16787
rect 15584 16772 15769 16786
rect 15584 16766 15587 16772
rect 15763 16770 15769 16772
rect 15786 16770 15792 16787
rect 15763 16767 15792 16770
rect 17073 16766 17076 16792
rect 17102 16766 17105 16792
rect 17257 16786 17260 16792
rect 17174 16772 17260 16786
rect 14635 16756 14638 16758
rect 14480 16753 14494 16756
rect 14488 16736 14494 16753
rect 14575 16753 14612 16756
rect 14480 16733 14494 16736
rect 14527 16748 14556 16751
rect 14480 16732 14483 16733
rect 14527 16731 14533 16748
rect 14550 16731 14556 16748
rect 14575 16736 14581 16753
rect 14598 16738 14612 16753
rect 14626 16753 14638 16756
rect 14598 16736 14604 16738
rect 14575 16733 14604 16736
rect 14626 16736 14632 16753
rect 14664 16752 14667 16758
rect 15509 16752 15512 16758
rect 14664 16738 15512 16752
rect 14626 16733 14638 16736
rect 14635 16732 14638 16733
rect 14664 16732 14667 16738
rect 15509 16732 15512 16738
rect 15538 16732 15541 16758
rect 15717 16753 15746 16756
rect 15717 16736 15723 16753
rect 15740 16752 15746 16753
rect 15831 16752 15834 16758
rect 15740 16738 15834 16752
rect 15740 16736 15746 16738
rect 15717 16733 15746 16736
rect 15831 16732 15834 16738
rect 15860 16732 15863 16758
rect 15969 16732 15972 16758
rect 15998 16752 16001 16758
rect 15998 16738 16544 16752
rect 15998 16732 16001 16738
rect 14527 16728 14556 16731
rect 14112 16704 14382 16718
rect 14112 16698 14115 16704
rect 8112 16670 9874 16684
rect 14532 16670 14546 16728
rect 15187 16698 15190 16724
rect 15216 16718 15219 16724
rect 15463 16718 15466 16724
rect 15216 16704 15466 16718
rect 15216 16698 15219 16704
rect 15463 16698 15466 16704
rect 15492 16718 15495 16724
rect 15556 16719 15585 16722
rect 15556 16718 15562 16719
rect 15492 16704 15562 16718
rect 15492 16698 15495 16704
rect 15556 16702 15562 16704
rect 15579 16702 15585 16719
rect 15556 16699 15585 16702
rect 16530 16690 16544 16738
rect 17119 16732 17122 16758
rect 17148 16752 17151 16758
rect 17174 16756 17188 16772
rect 17257 16766 17260 16772
rect 17286 16766 17289 16792
rect 17975 16787 18004 16790
rect 17975 16770 17981 16787
rect 17998 16786 18004 16787
rect 20229 16787 20258 16790
rect 17998 16772 18108 16786
rect 17998 16770 18004 16772
rect 17975 16767 18004 16770
rect 17166 16753 17195 16756
rect 17166 16752 17172 16753
rect 17148 16738 17172 16752
rect 17148 16732 17151 16738
rect 17166 16736 17172 16738
rect 17189 16736 17195 16753
rect 17166 16733 17195 16736
rect 17212 16753 17241 16756
rect 17212 16736 17218 16753
rect 17235 16736 17241 16753
rect 17212 16733 17241 16736
rect 17261 16748 17290 16751
rect 16591 16719 16620 16722
rect 16591 16702 16597 16719
rect 16614 16718 16620 16719
rect 17220 16718 17234 16733
rect 17261 16731 17267 16748
rect 17284 16731 17290 16748
rect 17717 16732 17720 16758
rect 17746 16752 17749 16758
rect 17764 16753 17793 16756
rect 17764 16752 17770 16753
rect 17746 16738 17770 16752
rect 17746 16732 17749 16738
rect 17764 16736 17770 16738
rect 17787 16736 17793 16753
rect 17764 16733 17793 16736
rect 17901 16732 17904 16758
rect 17930 16756 17933 16758
rect 17930 16753 17954 16756
rect 17930 16736 17931 16753
rect 17948 16736 17954 16753
rect 18094 16752 18108 16772
rect 20229 16770 20235 16787
rect 20252 16786 20258 16787
rect 21673 16786 21676 16792
rect 20252 16772 20362 16786
rect 20252 16770 20258 16772
rect 20109 16752 20112 16769
rect 18094 16743 20112 16752
rect 20138 16743 20141 16769
rect 20229 16767 20258 16770
rect 18094 16738 20132 16743
rect 17930 16733 17954 16736
rect 17930 16732 17933 16733
rect 20155 16732 20158 16758
rect 20184 16756 20187 16758
rect 20184 16753 20202 16756
rect 20196 16736 20202 16753
rect 20348 16752 20362 16772
rect 21575 16772 21676 16786
rect 20753 16752 20756 16758
rect 20348 16738 20756 16752
rect 20184 16733 20202 16736
rect 20184 16732 20187 16733
rect 20753 16732 20756 16738
rect 20782 16732 20785 16758
rect 21305 16732 21308 16758
rect 21334 16732 21337 16758
rect 21363 16753 21392 16756
rect 21363 16752 21369 16753
rect 21360 16736 21369 16752
rect 21386 16736 21392 16753
rect 21360 16733 21392 16736
rect 17261 16728 17290 16731
rect 16614 16704 17234 16718
rect 16614 16702 16620 16704
rect 16591 16699 16620 16702
rect 4745 16630 4748 16656
rect 4774 16650 4777 16656
rect 5021 16650 5024 16656
rect 4774 16636 5024 16650
rect 4774 16630 4777 16636
rect 5021 16630 5024 16636
rect 5050 16630 5053 16656
rect 6309 16630 6312 16656
rect 6338 16650 6341 16656
rect 8112 16650 8126 16670
rect 6338 16636 8126 16650
rect 8311 16651 8340 16654
rect 6338 16630 6341 16636
rect 8311 16634 8317 16651
rect 8334 16650 8340 16651
rect 8379 16650 8382 16656
rect 8334 16636 8382 16650
rect 8334 16634 8340 16636
rect 8311 16631 8340 16634
rect 8379 16630 8382 16636
rect 8408 16630 8411 16656
rect 9805 16630 9808 16656
rect 9834 16630 9837 16656
rect 9860 16650 9874 16670
rect 14543 16664 14546 16670
rect 14572 16664 14575 16690
rect 16521 16664 16524 16690
rect 16550 16684 16553 16690
rect 17266 16684 17280 16728
rect 20018 16719 20047 16722
rect 20018 16702 20024 16719
rect 20041 16702 20047 16719
rect 20018 16699 20047 16702
rect 21053 16719 21082 16722
rect 21053 16702 21059 16719
rect 21076 16718 21082 16719
rect 21360 16718 21374 16733
rect 21443 16732 21446 16758
rect 21472 16756 21475 16758
rect 21575 16756 21589 16772
rect 21673 16766 21676 16772
rect 21702 16766 21705 16792
rect 22915 16766 22918 16792
rect 22944 16786 22947 16792
rect 23169 16787 23198 16790
rect 23169 16786 23175 16787
rect 22944 16772 23175 16786
rect 22944 16766 22947 16772
rect 23169 16770 23175 16772
rect 23192 16770 23198 16787
rect 23169 16767 23198 16770
rect 25997 16766 26000 16792
rect 26026 16786 26029 16792
rect 26205 16787 26234 16790
rect 26205 16786 26211 16787
rect 26026 16772 26211 16786
rect 26026 16766 26029 16772
rect 26205 16770 26211 16772
rect 26228 16770 26234 16787
rect 26205 16767 26234 16770
rect 28343 16766 28346 16792
rect 28372 16786 28375 16792
rect 28550 16787 28579 16790
rect 28550 16786 28556 16787
rect 28372 16772 28556 16786
rect 28372 16766 28375 16772
rect 28550 16770 28556 16772
rect 28573 16770 28579 16787
rect 28550 16767 28579 16770
rect 28601 16787 28630 16790
rect 28601 16770 28607 16787
rect 28624 16786 28630 16787
rect 28665 16786 28668 16792
rect 28624 16772 28668 16786
rect 28624 16770 28630 16772
rect 28601 16767 28630 16770
rect 28665 16766 28668 16772
rect 28694 16766 28697 16792
rect 21472 16753 21486 16756
rect 21480 16736 21486 16753
rect 21567 16753 21596 16756
rect 21472 16733 21486 16736
rect 21519 16748 21548 16751
rect 21472 16732 21475 16733
rect 21519 16731 21525 16748
rect 21542 16731 21548 16748
rect 21567 16736 21573 16753
rect 21590 16736 21596 16753
rect 21567 16733 21596 16736
rect 21618 16753 21647 16756
rect 21618 16736 21624 16753
rect 21641 16752 21647 16753
rect 22685 16752 22688 16758
rect 21641 16738 22688 16752
rect 21641 16736 21647 16738
rect 21618 16733 21647 16736
rect 22685 16732 22688 16738
rect 22714 16732 22717 16758
rect 22777 16732 22780 16758
rect 22806 16752 22809 16758
rect 23099 16752 23102 16758
rect 23128 16756 23131 16758
rect 23128 16753 23146 16756
rect 22806 16738 23102 16752
rect 22806 16732 22809 16738
rect 23099 16732 23102 16738
rect 23140 16736 23146 16753
rect 23128 16733 23146 16736
rect 23128 16732 23131 16733
rect 26043 16732 26046 16758
rect 26072 16752 26075 16758
rect 26159 16753 26188 16756
rect 26159 16752 26165 16753
rect 26072 16738 26165 16752
rect 26072 16732 26075 16738
rect 26159 16736 26165 16738
rect 26182 16752 26188 16753
rect 26411 16752 26414 16758
rect 26182 16738 26414 16752
rect 26182 16736 26188 16738
rect 26159 16733 26188 16736
rect 26411 16732 26414 16738
rect 26440 16732 26443 16758
rect 28389 16732 28392 16758
rect 28418 16732 28421 16758
rect 21519 16728 21548 16731
rect 21076 16704 21374 16718
rect 21076 16702 21082 16704
rect 21053 16699 21082 16702
rect 16550 16670 17280 16684
rect 16550 16664 16553 16670
rect 11737 16650 11740 16656
rect 9860 16636 11740 16650
rect 11737 16630 11740 16636
rect 11766 16630 11769 16656
rect 12060 16651 12089 16654
rect 12060 16634 12066 16651
rect 12083 16650 12089 16651
rect 12151 16650 12154 16656
rect 12083 16636 12154 16650
rect 12083 16634 12089 16636
rect 12060 16631 12089 16634
rect 12151 16630 12154 16636
rect 12180 16630 12183 16656
rect 12795 16630 12798 16656
rect 12824 16650 12827 16656
rect 13025 16650 13028 16656
rect 12824 16636 13028 16650
rect 12824 16630 12827 16636
rect 13025 16630 13028 16636
rect 13054 16630 13057 16656
rect 15142 16651 15171 16654
rect 15142 16634 15148 16651
rect 15165 16650 15171 16651
rect 15877 16650 15880 16656
rect 15165 16636 15880 16650
rect 15165 16634 15171 16636
rect 15142 16631 15171 16634
rect 15877 16630 15880 16636
rect 15906 16630 15909 16656
rect 17074 16651 17103 16654
rect 17074 16634 17080 16651
rect 17097 16650 17103 16651
rect 17211 16650 17214 16656
rect 17097 16636 17214 16650
rect 17097 16634 17103 16636
rect 17074 16631 17103 16634
rect 17211 16630 17214 16636
rect 17240 16630 17243 16656
rect 20026 16650 20040 16699
rect 21527 16684 21541 16728
rect 22962 16719 22991 16722
rect 22962 16702 22968 16719
rect 22985 16702 22991 16719
rect 22962 16699 22991 16702
rect 25998 16719 26027 16722
rect 25998 16702 26004 16719
rect 26021 16702 26027 16719
rect 25998 16699 26027 16702
rect 21903 16684 21906 16690
rect 21527 16670 21906 16684
rect 21903 16664 21906 16670
rect 21932 16664 21935 16690
rect 20569 16650 20572 16656
rect 20026 16636 20572 16650
rect 20569 16630 20572 16636
rect 20598 16630 20601 16656
rect 22970 16650 22984 16699
rect 23145 16650 23148 16656
rect 22970 16636 23148 16650
rect 23145 16630 23148 16636
rect 23174 16630 23177 16656
rect 23997 16651 24026 16654
rect 23997 16634 24003 16651
rect 24020 16650 24026 16651
rect 24111 16650 24114 16656
rect 24020 16636 24114 16650
rect 24020 16634 24026 16636
rect 23997 16631 24026 16634
rect 24111 16630 24114 16636
rect 24140 16630 24143 16656
rect 26006 16650 26020 16699
rect 26687 16650 26690 16656
rect 26006 16636 26690 16650
rect 26687 16630 26690 16636
rect 26716 16630 26719 16656
rect 29425 16651 29454 16654
rect 29425 16634 29431 16651
rect 29448 16650 29454 16651
rect 29631 16650 29634 16656
rect 29448 16636 29634 16650
rect 29448 16634 29454 16636
rect 29425 16631 29454 16634
rect 29631 16630 29634 16636
rect 29660 16630 29663 16656
rect 3036 16568 29992 16616
rect 4745 16528 4748 16554
rect 4774 16548 4777 16554
rect 4774 16534 4860 16548
rect 4774 16528 4777 16534
rect 4654 16515 4683 16518
rect 4654 16498 4660 16515
rect 4677 16514 4683 16515
rect 4699 16514 4702 16520
rect 4677 16500 4702 16514
rect 4677 16498 4683 16500
rect 4654 16495 4683 16498
rect 4699 16494 4702 16500
rect 4728 16494 4731 16520
rect 4846 16480 4860 16534
rect 6769 16528 6772 16554
rect 6798 16548 6801 16554
rect 6798 16534 9483 16548
rect 6798 16528 6801 16534
rect 9469 16514 9483 16534
rect 9667 16528 9670 16554
rect 9696 16552 9699 16554
rect 9696 16549 9720 16552
rect 9696 16532 9697 16549
rect 9714 16532 9720 16549
rect 11623 16549 11652 16552
rect 9696 16529 9720 16532
rect 10320 16534 11576 16548
rect 9696 16528 9699 16529
rect 9469 16500 9667 16514
rect 4846 16466 4862 16480
rect 4653 16426 4656 16452
rect 4682 16426 4685 16452
rect 4745 16450 4748 16452
rect 4731 16447 4748 16450
rect 4731 16430 4737 16447
rect 4731 16427 4748 16430
rect 4745 16426 4748 16427
rect 4774 16426 4777 16452
rect 4848 16450 4862 16466
rect 4974 16466 5780 16480
rect 4805 16447 4834 16450
rect 4805 16446 4811 16447
rect 4800 16430 4811 16446
rect 4828 16430 4834 16447
rect 4848 16447 4882 16450
rect 4848 16432 4859 16447
rect 4800 16427 4834 16430
rect 4853 16430 4859 16432
rect 4876 16430 4882 16447
rect 4853 16427 4882 16430
rect 3687 16392 3690 16418
rect 3716 16412 3719 16418
rect 4561 16412 4564 16418
rect 3716 16398 4564 16412
rect 3716 16392 3719 16398
rect 4561 16392 4564 16398
rect 4590 16392 4593 16418
rect 4607 16392 4610 16418
rect 4636 16412 4639 16418
rect 4800 16412 4814 16427
rect 4914 16426 4917 16452
rect 4943 16426 4946 16452
rect 4974 16448 4988 16466
rect 4966 16445 4995 16448
rect 4966 16428 4972 16445
rect 4989 16428 4995 16445
rect 4966 16425 4995 16428
rect 5665 16426 5668 16452
rect 5694 16446 5697 16452
rect 5712 16447 5741 16450
rect 5712 16446 5718 16447
rect 5694 16432 5718 16446
rect 5694 16426 5697 16432
rect 5712 16430 5718 16432
rect 5735 16430 5741 16447
rect 5766 16446 5780 16466
rect 7275 16460 7278 16486
rect 7304 16480 7307 16486
rect 7644 16481 7673 16484
rect 7644 16480 7650 16481
rect 7304 16466 7650 16480
rect 7304 16460 7307 16466
rect 7644 16464 7650 16466
rect 7667 16464 7673 16481
rect 9653 16480 9667 16500
rect 9851 16494 9854 16520
rect 9880 16514 9883 16520
rect 10174 16515 10203 16518
rect 10174 16514 10180 16515
rect 9880 16500 10180 16514
rect 9880 16494 9883 16500
rect 10174 16498 10180 16500
rect 10197 16498 10203 16515
rect 10174 16495 10203 16498
rect 10320 16480 10334 16534
rect 11562 16514 11576 16534
rect 11623 16532 11629 16549
rect 11646 16548 11652 16549
rect 11691 16548 11694 16554
rect 11646 16534 11694 16548
rect 11646 16532 11652 16534
rect 11623 16529 11652 16532
rect 11691 16528 11694 16534
rect 11720 16528 11723 16554
rect 12473 16528 12476 16554
rect 12502 16548 12505 16554
rect 12502 16534 14704 16548
rect 12502 16528 12505 16534
rect 12243 16514 12246 16520
rect 11562 16500 12246 16514
rect 12243 16494 12246 16500
rect 12272 16494 12275 16520
rect 9653 16466 10334 16480
rect 7644 16461 7673 16464
rect 6309 16446 6312 16452
rect 5766 16432 6312 16446
rect 5712 16427 5741 16430
rect 6309 16426 6312 16432
rect 6338 16426 6341 16452
rect 7229 16426 7232 16452
rect 7258 16446 7261 16452
rect 7413 16446 7416 16452
rect 7258 16432 7416 16446
rect 7258 16426 7261 16432
rect 7413 16426 7416 16432
rect 7442 16426 7445 16452
rect 8012 16447 8041 16450
rect 8012 16430 8018 16447
rect 8035 16446 8041 16447
rect 8609 16446 8612 16452
rect 8035 16432 8612 16446
rect 8035 16430 8041 16432
rect 8012 16427 8041 16430
rect 8609 16426 8612 16432
rect 8638 16446 8641 16452
rect 8656 16447 8685 16450
rect 8656 16446 8662 16447
rect 8638 16432 8662 16446
rect 8638 16426 8641 16432
rect 8656 16430 8662 16432
rect 8679 16430 8685 16447
rect 8855 16447 8884 16450
rect 8855 16446 8861 16447
rect 8656 16427 8685 16430
rect 8756 16432 8861 16446
rect 4636 16398 4814 16412
rect 4636 16392 4639 16398
rect 5619 16392 5622 16418
rect 5648 16412 5651 16418
rect 5872 16413 5901 16416
rect 5872 16412 5878 16413
rect 5648 16398 5878 16412
rect 5648 16392 5651 16398
rect 5872 16396 5878 16398
rect 5895 16396 5901 16413
rect 5872 16393 5901 16396
rect 5923 16413 5952 16416
rect 5923 16396 5929 16413
rect 5946 16412 5952 16413
rect 5987 16412 5990 16418
rect 5946 16398 5990 16412
rect 5946 16396 5952 16398
rect 5923 16393 5952 16396
rect 5987 16392 5990 16398
rect 6016 16392 6019 16418
rect 7183 16392 7186 16418
rect 7212 16412 7215 16418
rect 8756 16412 8770 16432
rect 8855 16430 8861 16432
rect 8878 16446 8884 16447
rect 8878 16432 9690 16446
rect 8878 16430 8884 16432
rect 8855 16427 8884 16430
rect 7212 16398 8770 16412
rect 8816 16413 8845 16416
rect 7212 16392 7215 16398
rect 8816 16396 8822 16413
rect 8839 16412 8845 16413
rect 8931 16412 8934 16418
rect 8839 16398 8934 16412
rect 8839 16396 8845 16398
rect 8816 16393 8845 16396
rect 8931 16392 8934 16398
rect 8960 16392 8963 16418
rect 9676 16412 9690 16432
rect 9805 16426 9808 16452
rect 9834 16446 9837 16452
rect 10320 16450 10334 16466
rect 10587 16460 10590 16486
rect 10616 16460 10619 16486
rect 12749 16460 12752 16486
rect 12778 16480 12781 16486
rect 13808 16481 13837 16484
rect 13808 16480 13814 16481
rect 12778 16466 13814 16480
rect 12778 16460 12781 16466
rect 13808 16464 13814 16466
rect 13831 16464 13837 16481
rect 13808 16461 13837 16464
rect 10174 16447 10203 16450
rect 10174 16446 10180 16447
rect 9834 16432 10180 16446
rect 9834 16426 9837 16432
rect 10174 16430 10180 16432
rect 10197 16430 10203 16447
rect 10174 16427 10203 16430
rect 10312 16447 10341 16450
rect 10312 16430 10318 16447
rect 10335 16430 10341 16447
rect 10787 16447 10816 16450
rect 10787 16446 10793 16447
rect 10312 16427 10341 16430
rect 10366 16432 10793 16446
rect 10366 16412 10380 16432
rect 10787 16430 10793 16432
rect 10810 16446 10816 16447
rect 13163 16446 13166 16452
rect 10810 16432 13166 16446
rect 10810 16430 10816 16432
rect 10787 16427 10816 16430
rect 13163 16426 13166 16432
rect 13192 16426 13195 16452
rect 13945 16426 13948 16452
rect 13974 16450 13977 16452
rect 13974 16447 13992 16450
rect 13986 16430 13992 16447
rect 14497 16446 14500 16452
rect 13974 16427 13992 16430
rect 14138 16432 14500 16446
rect 13974 16426 13977 16427
rect 10748 16413 10777 16416
rect 10748 16412 10754 16413
rect 9676 16398 10380 16412
rect 10642 16398 10754 16412
rect 10642 16384 10656 16398
rect 10748 16396 10754 16398
rect 10771 16396 10777 16413
rect 10748 16393 10777 16396
rect 14019 16413 14048 16416
rect 14019 16396 14025 16413
rect 14042 16412 14048 16413
rect 14138 16412 14152 16432
rect 14497 16426 14500 16432
rect 14526 16426 14529 16452
rect 14690 16446 14704 16534
rect 14773 16528 14776 16554
rect 14802 16548 14805 16554
rect 14843 16549 14872 16552
rect 14843 16548 14849 16549
rect 14802 16534 14849 16548
rect 14802 16528 14805 16534
rect 14843 16532 14849 16534
rect 14866 16532 14872 16549
rect 14843 16529 14872 16532
rect 16959 16549 16988 16552
rect 16959 16532 16965 16549
rect 16982 16548 16988 16549
rect 17165 16548 17168 16554
rect 16982 16534 17168 16548
rect 16982 16532 16988 16534
rect 16959 16529 16988 16532
rect 17165 16528 17168 16534
rect 17194 16528 17197 16554
rect 20799 16528 20802 16554
rect 20828 16548 20831 16554
rect 22915 16548 22918 16554
rect 20828 16534 22918 16548
rect 20828 16528 20831 16534
rect 22915 16528 22918 16534
rect 22944 16528 22947 16554
rect 23974 16549 24003 16552
rect 23974 16532 23980 16549
rect 23997 16548 24003 16549
rect 24019 16548 24022 16554
rect 23997 16534 24022 16548
rect 23997 16532 24003 16534
rect 23974 16529 24003 16532
rect 24019 16528 24022 16534
rect 24048 16528 24051 16554
rect 29493 16528 29496 16554
rect 29522 16528 29525 16554
rect 22924 16514 22938 16528
rect 24709 16514 24712 16520
rect 22924 16500 24712 16514
rect 24709 16494 24712 16500
rect 24738 16514 24741 16520
rect 25583 16514 25586 16520
rect 24738 16500 25586 16514
rect 24738 16494 24741 16500
rect 25583 16494 25586 16500
rect 25612 16494 25615 16520
rect 15463 16460 15466 16486
rect 15492 16480 15495 16486
rect 15924 16481 15953 16484
rect 15924 16480 15930 16481
rect 15492 16466 15930 16480
rect 15492 16460 15495 16466
rect 15924 16464 15930 16466
rect 15947 16464 15953 16481
rect 15924 16461 15953 16464
rect 16079 16447 16108 16450
rect 16079 16446 16085 16447
rect 14690 16432 16085 16446
rect 15932 16418 15946 16432
rect 16079 16430 16085 16432
rect 16102 16430 16108 16447
rect 16079 16427 16108 16430
rect 16123 16447 16152 16450
rect 16123 16430 16129 16447
rect 16146 16446 16152 16447
rect 16199 16446 16202 16452
rect 16146 16432 16202 16446
rect 16146 16430 16152 16432
rect 16123 16427 16152 16430
rect 16199 16426 16202 16432
rect 16228 16426 16231 16452
rect 17211 16426 17214 16452
rect 17240 16426 17243 16452
rect 17303 16426 17306 16452
rect 17332 16426 17335 16452
rect 21305 16426 21308 16452
rect 21334 16446 21337 16452
rect 24066 16447 24095 16450
rect 24066 16446 24072 16447
rect 21334 16432 24072 16446
rect 21334 16426 21337 16432
rect 24066 16430 24072 16432
rect 24089 16430 24095 16447
rect 24066 16427 24095 16430
rect 14042 16398 14152 16412
rect 14042 16396 14048 16398
rect 14019 16393 14048 16396
rect 15923 16392 15926 16418
rect 15952 16392 15955 16418
rect 23973 16392 23976 16418
rect 24002 16392 24005 16418
rect 24074 16412 24088 16427
rect 24111 16426 24114 16452
rect 24140 16426 24143 16452
rect 24176 16447 24205 16450
rect 24176 16430 24182 16447
rect 24199 16446 24205 16447
rect 26089 16446 26092 16452
rect 24199 16432 26092 16446
rect 24199 16430 24205 16432
rect 24176 16427 24205 16430
rect 26089 16426 26092 16432
rect 26118 16426 26121 16452
rect 29585 16426 29588 16452
rect 29614 16426 29617 16452
rect 29631 16426 29634 16452
rect 29660 16426 29663 16452
rect 29677 16426 29680 16452
rect 29706 16450 29709 16452
rect 29706 16446 29710 16450
rect 29815 16446 29818 16452
rect 29706 16432 29818 16446
rect 29706 16427 29710 16432
rect 29706 16426 29709 16427
rect 29815 16426 29818 16432
rect 29844 16426 29847 16452
rect 25859 16412 25862 16418
rect 24074 16398 25862 16412
rect 25859 16392 25862 16398
rect 25888 16392 25891 16418
rect 29493 16392 29496 16418
rect 29522 16392 29525 16418
rect 6723 16358 6726 16384
rect 6752 16382 6755 16384
rect 6752 16379 6776 16382
rect 6752 16362 6753 16379
rect 6770 16362 6776 16379
rect 6752 16359 6776 16362
rect 6752 16358 6755 16359
rect 10265 16358 10268 16384
rect 10294 16358 10297 16384
rect 10633 16358 10636 16384
rect 10662 16358 10665 16384
rect 17257 16358 17260 16384
rect 17286 16358 17289 16384
rect 3036 16296 29992 16344
rect 4285 16280 4288 16282
rect 4263 16277 4288 16280
rect 4263 16260 4269 16277
rect 4286 16260 4288 16277
rect 4263 16257 4288 16260
rect 4285 16256 4288 16257
rect 4314 16256 4317 16282
rect 5021 16256 5024 16282
rect 5050 16276 5053 16282
rect 6402 16277 6431 16280
rect 5050 16262 6240 16276
rect 5050 16256 5053 16262
rect 4561 16222 4564 16248
rect 4590 16242 4593 16248
rect 6226 16246 6240 16262
rect 6402 16260 6408 16277
rect 6425 16276 6431 16277
rect 6425 16262 6654 16276
rect 6425 16260 6431 16262
rect 6402 16257 6431 16260
rect 6640 16246 6654 16262
rect 6723 16256 6726 16282
rect 6752 16256 6755 16282
rect 9829 16277 9858 16280
rect 9829 16260 9835 16277
rect 9852 16276 9858 16277
rect 10265 16276 10268 16282
rect 9852 16262 10268 16276
rect 9852 16260 9858 16262
rect 9829 16257 9858 16260
rect 10265 16256 10268 16262
rect 10294 16256 10297 16282
rect 13739 16277 13768 16280
rect 13739 16260 13745 16277
rect 13762 16276 13768 16277
rect 14451 16276 14454 16282
rect 13762 16262 14454 16276
rect 13762 16260 13768 16262
rect 13739 16257 13768 16260
rect 14451 16256 14454 16262
rect 14480 16256 14483 16282
rect 23859 16277 23888 16280
rect 23859 16260 23865 16277
rect 23882 16276 23888 16277
rect 23973 16276 23976 16282
rect 23882 16262 23976 16276
rect 23882 16260 23888 16262
rect 23859 16257 23888 16260
rect 23973 16256 23976 16262
rect 24002 16256 24005 16282
rect 29333 16277 29362 16280
rect 29333 16260 29339 16277
rect 29356 16276 29362 16277
rect 29493 16276 29496 16282
rect 29356 16262 29496 16276
rect 29356 16260 29362 16262
rect 29333 16257 29362 16260
rect 29493 16256 29496 16262
rect 29522 16256 29525 16282
rect 9023 16246 9026 16248
rect 4723 16243 4752 16246
rect 4723 16242 4729 16243
rect 4590 16228 4729 16242
rect 4590 16222 4593 16228
rect 4723 16226 4729 16228
rect 4746 16226 4752 16243
rect 4723 16223 4752 16226
rect 6218 16243 6247 16246
rect 6218 16226 6224 16243
rect 6241 16226 6247 16243
rect 6218 16223 6247 16226
rect 6632 16243 6661 16246
rect 6632 16226 6638 16243
rect 6655 16226 6661 16243
rect 6632 16223 6661 16226
rect 7441 16243 7470 16246
rect 7441 16226 7447 16243
rect 7464 16242 7470 16243
rect 9005 16243 9026 16246
rect 7464 16228 7574 16242
rect 7464 16226 7470 16228
rect 7441 16223 7470 16226
rect 3135 16188 3138 16214
rect 3164 16208 3167 16214
rect 3228 16209 3257 16212
rect 3228 16208 3234 16209
rect 3164 16194 3234 16208
rect 3164 16188 3167 16194
rect 3228 16192 3234 16194
rect 3251 16192 3257 16209
rect 3228 16189 3257 16192
rect 3365 16188 3368 16214
rect 3394 16212 3397 16214
rect 3394 16209 3412 16212
rect 3406 16192 3412 16209
rect 3394 16189 3412 16192
rect 3427 16209 3456 16212
rect 3427 16192 3433 16209
rect 3450 16208 3456 16209
rect 4469 16208 4472 16214
rect 3450 16194 4472 16208
rect 3450 16192 3456 16194
rect 3427 16189 3456 16192
rect 3394 16188 3397 16189
rect 4469 16188 4472 16194
rect 4498 16188 4501 16214
rect 4515 16188 4518 16214
rect 4544 16188 4547 16214
rect 4677 16209 4706 16212
rect 4677 16192 4683 16209
rect 4700 16208 4706 16209
rect 4791 16208 4794 16214
rect 4700 16194 4794 16208
rect 4700 16192 4706 16194
rect 4677 16189 4706 16192
rect 4791 16188 4794 16194
rect 4820 16188 4823 16214
rect 5551 16209 5580 16212
rect 5551 16192 5557 16209
rect 5574 16208 5580 16209
rect 6126 16209 6155 16212
rect 6126 16208 6132 16209
rect 5574 16194 6132 16208
rect 5574 16192 5580 16194
rect 5551 16189 5580 16192
rect 6126 16192 6132 16194
rect 6149 16192 6155 16209
rect 6126 16189 6155 16192
rect 6263 16188 6266 16214
rect 6292 16188 6295 16214
rect 6309 16188 6312 16214
rect 6338 16188 6341 16214
rect 6769 16188 6772 16214
rect 6798 16188 6801 16214
rect 7230 16209 7259 16212
rect 7230 16192 7236 16209
rect 7253 16208 7259 16209
rect 7275 16208 7278 16214
rect 7253 16194 7278 16208
rect 7253 16192 7259 16194
rect 7230 16189 7259 16192
rect 7275 16188 7278 16194
rect 7304 16188 7307 16214
rect 7391 16209 7420 16212
rect 7391 16192 7397 16209
rect 7414 16208 7420 16209
rect 7505 16208 7508 16214
rect 7414 16194 7508 16208
rect 7414 16192 7420 16194
rect 7391 16189 7420 16192
rect 7505 16188 7508 16194
rect 7534 16188 7537 16214
rect 7560 16208 7574 16228
rect 9005 16226 9011 16243
rect 9005 16223 9026 16226
rect 9023 16222 9026 16223
rect 9052 16222 9055 16248
rect 12933 16246 12936 16248
rect 12915 16243 12936 16246
rect 12915 16226 12921 16243
rect 12915 16223 12936 16226
rect 12933 16222 12936 16223
rect 12962 16222 12965 16248
rect 20799 16222 20802 16248
rect 20828 16242 20831 16248
rect 20961 16243 20990 16246
rect 20961 16242 20967 16243
rect 20828 16228 20967 16242
rect 20828 16222 20831 16228
rect 20961 16226 20967 16228
rect 20984 16226 20990 16243
rect 23035 16243 23064 16246
rect 23035 16242 23041 16243
rect 20961 16223 20990 16226
rect 21774 16228 23041 16242
rect 8241 16208 8244 16214
rect 7560 16194 8244 16208
rect 8241 16188 8244 16194
rect 8270 16208 8273 16214
rect 8471 16208 8474 16214
rect 8270 16194 8474 16208
rect 8270 16188 8273 16194
rect 8471 16188 8474 16194
rect 8500 16188 8503 16214
rect 8609 16188 8612 16214
rect 8638 16208 8641 16214
rect 8794 16209 8823 16212
rect 8794 16208 8800 16209
rect 8638 16194 8800 16208
rect 8638 16188 8641 16194
rect 8794 16192 8800 16194
rect 8817 16192 8823 16209
rect 8794 16189 8823 16192
rect 8931 16188 8934 16214
rect 8960 16212 8963 16214
rect 8960 16209 8978 16212
rect 8972 16192 8978 16209
rect 8960 16189 8978 16192
rect 12704 16209 12733 16212
rect 12704 16192 12710 16209
rect 12727 16208 12733 16209
rect 12749 16208 12752 16214
rect 12727 16194 12752 16208
rect 12727 16192 12733 16194
rect 12704 16189 12733 16192
rect 8960 16188 8963 16189
rect 12749 16188 12752 16194
rect 12778 16188 12781 16214
rect 12841 16188 12844 16214
rect 12870 16212 12873 16214
rect 12870 16209 12888 16212
rect 12882 16192 12888 16209
rect 12870 16189 12888 16192
rect 20915 16209 20944 16212
rect 20915 16192 20921 16209
rect 20938 16208 20944 16209
rect 21029 16208 21032 16214
rect 20938 16194 21032 16208
rect 20938 16192 20944 16194
rect 20915 16189 20944 16192
rect 12870 16188 12873 16189
rect 21029 16188 21032 16194
rect 21058 16188 21061 16214
rect 20569 16154 20572 16180
rect 20598 16174 20601 16180
rect 20754 16175 20783 16178
rect 20754 16174 20760 16175
rect 20598 16160 20760 16174
rect 20598 16154 20601 16160
rect 20754 16158 20760 16160
rect 20777 16158 20783 16175
rect 20754 16155 20783 16158
rect 7183 16140 7186 16146
rect 5398 16126 7186 16140
rect 5398 16112 5412 16126
rect 7183 16120 7186 16126
rect 7212 16120 7215 16146
rect 21774 16140 21788 16228
rect 23035 16226 23041 16228
rect 23058 16242 23064 16243
rect 23058 16226 23076 16242
rect 23035 16223 23076 16226
rect 22777 16188 22780 16214
rect 22806 16208 22809 16214
rect 22979 16209 23008 16212
rect 22979 16208 22985 16209
rect 22806 16194 22985 16208
rect 22806 16188 22809 16194
rect 22979 16192 22985 16194
rect 23002 16192 23008 16209
rect 23062 16208 23076 16223
rect 25905 16222 25908 16248
rect 25934 16242 25937 16248
rect 26113 16243 26142 16246
rect 26113 16242 26119 16243
rect 25934 16228 26119 16242
rect 25934 16222 25937 16228
rect 26113 16226 26119 16228
rect 26136 16226 26142 16243
rect 26113 16223 26142 16226
rect 28297 16222 28300 16248
rect 28326 16242 28329 16248
rect 28505 16243 28534 16246
rect 28505 16242 28511 16243
rect 28326 16228 28511 16242
rect 28326 16222 28329 16228
rect 28505 16226 28511 16228
rect 28528 16226 28534 16243
rect 28505 16223 28534 16226
rect 24525 16208 24528 16214
rect 23062 16194 24528 16208
rect 22979 16189 23008 16192
rect 24525 16188 24528 16194
rect 24554 16188 24557 16214
rect 26043 16188 26046 16214
rect 26072 16212 26075 16214
rect 26072 16209 26090 16212
rect 26084 16192 26090 16209
rect 26072 16189 26090 16192
rect 26072 16188 26075 16189
rect 28343 16188 28346 16214
rect 28372 16208 28375 16214
rect 28453 16209 28482 16212
rect 28453 16208 28459 16209
rect 28372 16194 28459 16208
rect 28372 16188 28375 16194
rect 28453 16192 28459 16194
rect 28476 16192 28482 16209
rect 28453 16189 28482 16192
rect 22824 16175 22853 16178
rect 22824 16158 22830 16175
rect 22847 16158 22853 16175
rect 22824 16155 22853 16158
rect 21590 16126 21788 16140
rect 4515 16086 4518 16112
rect 4544 16106 4547 16112
rect 5389 16106 5392 16112
rect 4544 16092 5392 16106
rect 4544 16086 4547 16092
rect 5389 16086 5392 16092
rect 5418 16086 5421 16112
rect 6631 16086 6634 16112
rect 6660 16086 6663 16112
rect 8195 16086 8198 16112
rect 8224 16106 8227 16112
rect 8265 16107 8294 16110
rect 8265 16106 8271 16107
rect 8224 16092 8271 16106
rect 8224 16086 8227 16092
rect 8265 16090 8271 16092
rect 8288 16090 8294 16107
rect 8265 16087 8294 16090
rect 20753 16086 20756 16112
rect 20782 16106 20785 16112
rect 21590 16106 21604 16126
rect 20782 16092 21604 16106
rect 21789 16107 21818 16110
rect 20782 16086 20785 16092
rect 21789 16090 21795 16107
rect 21812 16106 21818 16107
rect 21857 16106 21860 16112
rect 21812 16092 21860 16106
rect 21812 16090 21818 16092
rect 21789 16087 21818 16090
rect 21857 16086 21860 16092
rect 21886 16086 21889 16112
rect 22832 16106 22846 16155
rect 25353 16154 25356 16180
rect 25382 16174 25385 16180
rect 25906 16175 25935 16178
rect 25906 16174 25912 16175
rect 25382 16160 25912 16174
rect 25382 16154 25385 16160
rect 25906 16158 25912 16160
rect 25929 16158 25935 16175
rect 25906 16155 25935 16158
rect 23145 16106 23148 16112
rect 22832 16092 23148 16106
rect 23145 16086 23148 16092
rect 23174 16086 23177 16112
rect 25914 16106 25928 16155
rect 28297 16154 28300 16180
rect 28326 16154 28329 16180
rect 26733 16106 26736 16112
rect 25914 16092 26736 16106
rect 26733 16086 26736 16092
rect 26762 16086 26765 16112
rect 26941 16107 26970 16110
rect 26941 16090 26947 16107
rect 26964 16106 26970 16107
rect 27193 16106 27196 16112
rect 26964 16092 27196 16106
rect 26964 16090 26970 16092
rect 26941 16087 26970 16090
rect 27193 16086 27196 16092
rect 27222 16086 27225 16112
rect 3036 16024 29992 16072
rect 4171 16005 4200 16008
rect 4171 15988 4177 16005
rect 4194 16004 4200 16005
rect 4653 16004 4656 16010
rect 4194 15990 4656 16004
rect 4194 15988 4200 15990
rect 4171 15985 4200 15988
rect 4653 15984 4656 15990
rect 4682 15984 4685 16010
rect 6195 16005 6224 16008
rect 6195 15988 6201 16005
rect 6218 16004 6224 16005
rect 6263 16004 6266 16010
rect 6218 15990 6266 16004
rect 6218 15988 6224 15990
rect 6195 15985 6224 15988
rect 6263 15984 6266 15990
rect 6292 15984 6295 16010
rect 8977 16004 8980 16010
rect 8112 15990 8980 16004
rect 3135 15916 3138 15942
rect 3164 15916 3167 15942
rect 3297 15903 3326 15906
rect 3297 15886 3303 15903
rect 3320 15902 3326 15903
rect 3411 15902 3414 15908
rect 3320 15888 3414 15902
rect 3320 15886 3326 15888
rect 3297 15883 3326 15886
rect 3411 15882 3414 15888
rect 3440 15882 3443 15908
rect 4791 15882 4794 15908
rect 4820 15902 4823 15908
rect 5160 15903 5189 15906
rect 4820 15882 4837 15902
rect 5160 15886 5166 15903
rect 5183 15902 5189 15903
rect 5711 15902 5714 15908
rect 5183 15888 5714 15902
rect 5183 15886 5189 15888
rect 5160 15883 5189 15886
rect 5711 15882 5714 15888
rect 5740 15882 5743 15908
rect 5757 15882 5760 15908
rect 5786 15902 5789 15908
rect 7505 15902 7508 15908
rect 5786 15888 7508 15902
rect 5786 15882 5789 15888
rect 7505 15882 7508 15888
rect 7534 15882 7537 15908
rect 8112 15906 8126 15990
rect 8977 15984 8980 15990
rect 9006 16004 9009 16010
rect 9299 16004 9302 16010
rect 9006 15990 9302 16004
rect 9006 15984 9009 15990
rect 9299 15984 9302 15990
rect 9328 15984 9331 16010
rect 8287 15950 8290 15976
rect 8316 15950 8319 15976
rect 25813 15950 25816 15976
rect 25842 15970 25845 15976
rect 25842 15956 25974 15970
rect 25842 15950 25845 15956
rect 8296 15936 8310 15950
rect 8250 15922 8310 15936
rect 10688 15922 10840 15936
rect 8195 15906 8198 15908
rect 8104 15903 8133 15906
rect 8104 15886 8110 15903
rect 8127 15886 8133 15903
rect 8104 15883 8133 15886
rect 8181 15903 8198 15906
rect 8181 15886 8187 15903
rect 8181 15883 8198 15886
rect 8195 15882 8198 15883
rect 8224 15882 8227 15908
rect 8250 15904 8264 15922
rect 8250 15901 8284 15904
rect 8250 15888 8261 15901
rect 8255 15884 8261 15888
rect 8278 15884 8284 15901
rect 8365 15903 8394 15906
rect 3365 15872 3368 15874
rect 3347 15869 3368 15872
rect 3347 15852 3353 15869
rect 3347 15849 3368 15852
rect 3365 15848 3368 15849
rect 3394 15848 3397 15874
rect 4823 15868 4837 15882
rect 8255 15881 8284 15884
rect 8311 15893 8340 15896
rect 8311 15876 8317 15893
rect 8334 15876 8340 15893
rect 8365 15886 8371 15903
rect 8388 15902 8394 15903
rect 8416 15903 8445 15906
rect 8388 15886 8402 15902
rect 8365 15883 8402 15886
rect 8416 15886 8422 15903
rect 8439 15902 8445 15903
rect 9207 15902 9210 15908
rect 8439 15888 9210 15902
rect 8439 15886 8445 15888
rect 8416 15883 8445 15886
rect 5205 15868 5208 15874
rect 4823 15854 5208 15868
rect 5205 15848 5208 15854
rect 5234 15868 5237 15874
rect 5389 15872 5392 15874
rect 5320 15869 5349 15872
rect 5320 15868 5326 15869
rect 5234 15854 5326 15868
rect 5234 15848 5237 15854
rect 5320 15852 5326 15854
rect 5343 15852 5349 15869
rect 5320 15849 5349 15852
rect 5371 15869 5392 15872
rect 5371 15852 5377 15869
rect 5371 15849 5392 15852
rect 5389 15848 5392 15849
rect 5418 15848 5421 15874
rect 8311 15873 8340 15876
rect 8319 15840 8333 15873
rect 8388 15840 8402 15883
rect 9207 15882 9210 15888
rect 9236 15882 9239 15908
rect 9345 15848 9348 15874
rect 9374 15868 9377 15874
rect 10688 15868 10702 15922
rect 10771 15882 10774 15908
rect 10800 15882 10803 15908
rect 10826 15902 10840 15922
rect 25353 15916 25356 15942
rect 25382 15916 25385 15942
rect 25583 15916 25586 15942
rect 25612 15936 25615 15942
rect 25859 15936 25862 15942
rect 25612 15922 25862 15936
rect 25612 15916 25615 15922
rect 25853 15916 25862 15922
rect 25888 15916 25891 15942
rect 25960 15936 25974 15956
rect 26089 15936 26092 15942
rect 25960 15922 26092 15936
rect 10971 15903 11000 15906
rect 10971 15902 10977 15903
rect 10826 15888 10977 15902
rect 10971 15886 10977 15888
rect 10994 15886 11000 15903
rect 10971 15883 11000 15886
rect 24157 15882 24160 15908
rect 24186 15902 24189 15908
rect 24342 15903 24371 15906
rect 24342 15902 24348 15903
rect 24186 15888 24348 15902
rect 24186 15882 24189 15888
rect 24342 15886 24348 15888
rect 24365 15902 24371 15903
rect 25362 15902 25376 15916
rect 24365 15888 25376 15902
rect 24365 15886 24371 15888
rect 24342 15883 24371 15886
rect 25629 15882 25632 15908
rect 25658 15882 25661 15908
rect 25721 15906 25724 15908
rect 25707 15903 25724 15906
rect 25707 15886 25713 15903
rect 25707 15883 25724 15886
rect 25721 15882 25724 15883
rect 25750 15882 25753 15908
rect 25788 15903 25817 15906
rect 25788 15886 25794 15903
rect 25811 15886 25817 15903
rect 25853 15896 25867 15916
rect 25960 15906 25974 15922
rect 26089 15916 26092 15922
rect 26118 15916 26121 15942
rect 26733 15916 26736 15942
rect 26762 15916 26765 15942
rect 29309 15936 29312 15942
rect 28720 15922 29312 15936
rect 25942 15903 25974 15906
rect 25788 15883 25817 15886
rect 25843 15893 25872 15896
rect 9374 15854 10702 15868
rect 9374 15848 9377 15854
rect 10817 15848 10820 15874
rect 10846 15868 10849 15874
rect 10932 15869 10961 15872
rect 10932 15868 10938 15869
rect 10846 15854 10938 15868
rect 10846 15848 10849 15854
rect 10932 15852 10938 15854
rect 10955 15852 10961 15869
rect 10932 15849 10961 15852
rect 24387 15848 24390 15874
rect 24416 15868 24419 15874
rect 24571 15872 24574 15874
rect 24502 15869 24531 15872
rect 24502 15868 24508 15869
rect 24416 15854 24508 15868
rect 24416 15848 24419 15854
rect 24502 15852 24508 15854
rect 24525 15852 24531 15869
rect 24502 15849 24531 15852
rect 24553 15869 24574 15872
rect 24553 15852 24559 15869
rect 24553 15849 24574 15852
rect 24571 15848 24574 15849
rect 24600 15848 24603 15874
rect 25377 15869 25406 15872
rect 25377 15852 25383 15869
rect 25400 15868 25406 15869
rect 25789 15868 25803 15883
rect 25843 15876 25849 15893
rect 25866 15876 25872 15893
rect 25843 15873 25872 15876
rect 25891 15893 25920 15896
rect 25891 15876 25897 15893
rect 25914 15891 25920 15893
rect 25914 15876 25928 15891
rect 25942 15886 25948 15903
rect 25965 15888 25974 15903
rect 26365 15902 26368 15908
rect 26006 15888 26368 15902
rect 25965 15886 25971 15888
rect 25942 15883 25971 15886
rect 25891 15873 25928 15876
rect 25400 15854 25803 15868
rect 25914 15868 25928 15873
rect 26006 15868 26020 15888
rect 26365 15882 26368 15888
rect 26394 15882 26397 15908
rect 28159 15882 28162 15908
rect 28188 15902 28191 15908
rect 28720 15906 28734 15922
rect 29309 15916 29312 15922
rect 29338 15916 29341 15942
rect 28712 15903 28741 15906
rect 28188 15888 28688 15902
rect 28188 15882 28191 15888
rect 25914 15854 26020 15868
rect 25400 15852 25406 15854
rect 25377 15849 25406 15852
rect 26043 15848 26046 15874
rect 26072 15868 26075 15874
rect 26779 15868 26782 15874
rect 26072 15854 26782 15868
rect 26072 15848 26075 15854
rect 26779 15848 26782 15854
rect 26808 15868 26811 15874
rect 26895 15869 26924 15872
rect 26895 15868 26901 15869
rect 26808 15854 26901 15868
rect 26808 15848 26811 15854
rect 26895 15852 26901 15854
rect 26918 15852 26924 15869
rect 26895 15849 26924 15852
rect 26945 15869 26974 15872
rect 26945 15852 26951 15869
rect 26968 15868 26974 15869
rect 27009 15868 27012 15874
rect 26968 15854 27012 15868
rect 26968 15852 26974 15854
rect 26945 15849 26974 15852
rect 27009 15848 27012 15854
rect 27038 15848 27041 15874
rect 7229 15814 7232 15840
rect 7258 15834 7261 15840
rect 8104 15835 8133 15838
rect 8104 15834 8110 15835
rect 7258 15820 8110 15834
rect 7258 15814 7261 15820
rect 8104 15818 8110 15820
rect 8127 15818 8133 15835
rect 8104 15815 8133 15818
rect 8241 15814 8244 15840
rect 8270 15834 8273 15840
rect 8319 15834 8336 15840
rect 8270 15820 8336 15834
rect 8270 15814 8273 15820
rect 8333 15814 8336 15820
rect 8362 15814 8365 15840
rect 8379 15814 8382 15840
rect 8408 15814 8411 15840
rect 10633 15814 10636 15840
rect 10662 15834 10665 15840
rect 10826 15834 10840 15848
rect 11829 15838 11832 15840
rect 10662 15820 10840 15834
rect 11807 15835 11832 15838
rect 10662 15814 10665 15820
rect 11807 15818 11813 15835
rect 11830 15818 11832 15835
rect 11807 15815 11832 15818
rect 11829 15814 11832 15815
rect 11858 15814 11861 15840
rect 20983 15814 20986 15840
rect 21012 15834 21015 15840
rect 22961 15834 22964 15840
rect 21012 15820 22964 15834
rect 21012 15814 21015 15820
rect 22961 15814 22964 15820
rect 22990 15814 22993 15840
rect 25860 15835 25889 15838
rect 25860 15818 25866 15835
rect 25883 15834 25889 15835
rect 26503 15834 26506 15840
rect 25883 15820 26506 15834
rect 25883 15818 25889 15820
rect 25860 15815 25889 15818
rect 26503 15814 26506 15820
rect 26532 15814 26535 15840
rect 27285 15814 27288 15840
rect 27314 15834 27317 15840
rect 27769 15835 27798 15838
rect 27769 15834 27775 15835
rect 27314 15820 27775 15834
rect 27314 15814 27317 15820
rect 27769 15818 27775 15820
rect 27792 15818 27798 15835
rect 28674 15834 28688 15888
rect 28712 15886 28718 15903
rect 28735 15886 28741 15903
rect 28712 15883 28741 15886
rect 28804 15903 28833 15906
rect 28804 15886 28810 15903
rect 28827 15886 28833 15903
rect 28804 15883 28833 15886
rect 28942 15903 28971 15906
rect 28942 15886 28948 15903
rect 28965 15902 28971 15903
rect 28987 15902 28990 15908
rect 28965 15888 28990 15902
rect 28965 15886 28971 15888
rect 28942 15883 28971 15886
rect 28757 15848 28760 15874
rect 28786 15848 28789 15874
rect 28812 15834 28826 15883
rect 28987 15882 28990 15888
rect 29016 15882 29019 15908
rect 28674 15820 28826 15834
rect 27769 15815 27798 15818
rect 3036 15752 29992 15800
rect 4493 15733 4522 15736
rect 4493 15716 4499 15733
rect 4516 15732 4522 15733
rect 4607 15732 4610 15738
rect 4516 15718 4610 15732
rect 4516 15716 4522 15718
rect 4493 15713 4522 15716
rect 4607 15712 4610 15718
rect 4636 15712 4639 15738
rect 5205 15712 5208 15738
rect 5234 15732 5237 15738
rect 5619 15732 5622 15738
rect 5234 15718 5622 15732
rect 5234 15712 5237 15718
rect 5619 15712 5622 15718
rect 5648 15712 5651 15738
rect 21857 15732 21860 15738
rect 21851 15712 21860 15732
rect 21886 15712 21889 15738
rect 26365 15712 26368 15738
rect 26394 15736 26397 15738
rect 26394 15733 26418 15736
rect 26394 15716 26395 15733
rect 26412 15716 26418 15733
rect 26394 15713 26418 15716
rect 27378 15733 27407 15736
rect 27378 15716 27384 15733
rect 27401 15732 27407 15733
rect 28159 15732 28162 15738
rect 27401 15718 28162 15732
rect 27401 15716 27407 15718
rect 27378 15713 27407 15716
rect 26394 15712 26397 15713
rect 28159 15712 28162 15718
rect 28188 15712 28191 15738
rect 3687 15702 3690 15704
rect 3669 15699 3690 15702
rect 3669 15682 3675 15699
rect 3669 15679 3690 15682
rect 3687 15678 3690 15679
rect 3716 15678 3719 15704
rect 8425 15678 8428 15704
rect 8454 15698 8457 15704
rect 9419 15699 9448 15702
rect 9419 15698 9425 15699
rect 8454 15684 9425 15698
rect 8454 15678 8457 15684
rect 9419 15682 9425 15684
rect 9442 15698 9448 15699
rect 11093 15698 11096 15704
rect 9442 15682 9460 15698
rect 9419 15679 9460 15682
rect 3411 15644 3414 15670
rect 3440 15664 3443 15670
rect 3619 15665 3648 15668
rect 3619 15664 3625 15665
rect 3440 15650 3625 15664
rect 3440 15644 3443 15650
rect 3619 15648 3625 15650
rect 3642 15664 3648 15665
rect 5665 15664 5668 15670
rect 3642 15650 5668 15664
rect 3642 15648 3648 15650
rect 3619 15645 3648 15648
rect 5665 15644 5668 15650
rect 5694 15664 5697 15670
rect 5757 15664 5760 15670
rect 5694 15650 5760 15664
rect 5694 15644 5697 15650
rect 5757 15644 5760 15650
rect 5786 15644 5789 15670
rect 9023 15644 9026 15670
rect 9052 15664 9055 15670
rect 9253 15664 9256 15670
rect 9052 15650 9256 15664
rect 9052 15644 9055 15650
rect 9253 15644 9256 15650
rect 9282 15664 9285 15670
rect 9363 15665 9392 15668
rect 9363 15664 9369 15665
rect 9282 15650 9369 15664
rect 9282 15644 9285 15650
rect 9363 15648 9369 15650
rect 9386 15648 9392 15665
rect 9446 15664 9460 15679
rect 11033 15684 11096 15698
rect 11033 15664 11047 15684
rect 11093 15678 11096 15684
rect 11122 15698 11125 15704
rect 12685 15699 12714 15702
rect 12685 15698 12691 15699
rect 11122 15684 12691 15698
rect 11122 15678 11125 15684
rect 12685 15682 12691 15684
rect 12708 15698 12714 15699
rect 12708 15682 12726 15698
rect 12685 15679 12726 15682
rect 9446 15650 11047 15664
rect 9363 15645 9392 15648
rect 12519 15644 12522 15670
rect 12548 15664 12551 15670
rect 12629 15665 12658 15668
rect 12629 15664 12635 15665
rect 12548 15650 12635 15664
rect 12548 15644 12551 15650
rect 12629 15648 12635 15650
rect 12652 15648 12658 15665
rect 12712 15664 12726 15679
rect 15371 15678 15374 15704
rect 15400 15698 15403 15704
rect 18527 15699 18556 15702
rect 15400 15684 15546 15698
rect 15400 15678 15403 15684
rect 13025 15664 13028 15670
rect 12712 15650 13028 15664
rect 12629 15645 12658 15648
rect 13025 15644 13028 15650
rect 13054 15644 13057 15670
rect 15463 15644 15466 15670
rect 15492 15668 15495 15670
rect 15532 15668 15546 15684
rect 18527 15682 18533 15699
rect 18550 15698 18556 15699
rect 18591 15698 18594 15704
rect 18550 15684 18594 15698
rect 18550 15682 18556 15684
rect 18527 15679 18556 15682
rect 18591 15678 18594 15684
rect 18620 15678 18623 15704
rect 20109 15678 20112 15704
rect 20138 15698 20141 15704
rect 20293 15702 20296 15704
rect 20275 15699 20296 15702
rect 20275 15698 20281 15699
rect 20138 15684 20281 15698
rect 20138 15678 20141 15684
rect 20275 15682 20281 15684
rect 20275 15679 20296 15682
rect 20293 15678 20296 15679
rect 20322 15678 20325 15704
rect 21851 15679 21865 15712
rect 21843 15676 21872 15679
rect 24387 15678 24390 15704
rect 24416 15698 24419 15704
rect 25583 15702 25586 15704
rect 25565 15699 25586 15702
rect 24416 15684 25537 15698
rect 24416 15678 24419 15684
rect 15492 15665 15510 15668
rect 15504 15648 15510 15665
rect 15492 15645 15510 15648
rect 15525 15665 15554 15668
rect 15525 15648 15531 15665
rect 15548 15664 15554 15665
rect 16199 15664 16202 15670
rect 15548 15650 16202 15664
rect 15548 15648 15554 15650
rect 15525 15645 15554 15648
rect 15492 15644 15495 15645
rect 16199 15644 16202 15650
rect 16228 15644 16231 15670
rect 18477 15665 18506 15668
rect 18477 15648 18483 15665
rect 18500 15664 18506 15665
rect 18729 15664 18732 15670
rect 18500 15650 18732 15664
rect 18500 15648 18506 15650
rect 18477 15645 18506 15648
rect 18729 15644 18732 15650
rect 18758 15664 18761 15670
rect 20225 15665 20254 15668
rect 20225 15664 20231 15665
rect 18758 15650 20231 15664
rect 18758 15644 18761 15650
rect 20225 15648 20231 15650
rect 20248 15664 20254 15665
rect 20799 15664 20802 15670
rect 20248 15650 20802 15664
rect 20248 15648 20254 15650
rect 20225 15645 20254 15648
rect 20799 15644 20802 15650
rect 20828 15664 20831 15670
rect 21099 15665 21128 15668
rect 20828 15650 21052 15664
rect 20828 15644 20831 15650
rect 21038 15636 21052 15650
rect 21099 15648 21105 15665
rect 21122 15664 21128 15665
rect 21582 15665 21611 15668
rect 21582 15664 21588 15665
rect 21122 15650 21588 15664
rect 21122 15648 21128 15650
rect 21099 15645 21128 15648
rect 21582 15648 21588 15650
rect 21605 15648 21611 15665
rect 21582 15645 21611 15648
rect 21627 15644 21630 15670
rect 21656 15668 21659 15670
rect 21656 15665 21668 15668
rect 21662 15648 21668 15665
rect 21656 15645 21668 15648
rect 21656 15644 21659 15645
rect 21719 15644 21722 15670
rect 21748 15668 21751 15670
rect 21748 15665 21762 15668
rect 21756 15648 21762 15665
rect 21748 15645 21762 15648
rect 21789 15665 21818 15668
rect 21789 15648 21795 15665
rect 21812 15648 21818 15665
rect 21843 15659 21849 15676
rect 21866 15659 21872 15676
rect 21903 15668 21906 15670
rect 21843 15656 21872 15659
rect 21894 15665 21906 15668
rect 21789 15645 21818 15648
rect 21894 15648 21900 15665
rect 21894 15645 21906 15648
rect 21748 15644 21751 15645
rect 3135 15610 3138 15636
rect 3164 15630 3167 15636
rect 3457 15630 3460 15636
rect 3164 15616 3460 15630
rect 3164 15610 3167 15616
rect 3457 15610 3460 15616
rect 3486 15610 3489 15636
rect 9115 15610 9118 15636
rect 9144 15630 9147 15636
rect 9208 15631 9237 15634
rect 9208 15630 9214 15631
rect 9144 15616 9214 15630
rect 9144 15610 9147 15616
rect 9208 15614 9214 15616
rect 9231 15614 9237 15631
rect 9208 15611 9237 15614
rect 12381 15610 12384 15636
rect 12410 15630 12413 15636
rect 12474 15631 12503 15634
rect 12474 15630 12480 15631
rect 12410 15616 12480 15630
rect 12410 15610 12413 15616
rect 12474 15614 12480 15616
rect 12497 15614 12503 15631
rect 12474 15611 12503 15614
rect 15187 15610 15190 15636
rect 15216 15630 15219 15636
rect 15326 15631 15355 15634
rect 15326 15630 15332 15631
rect 15216 15616 15332 15630
rect 15216 15610 15219 15616
rect 15326 15614 15332 15616
rect 15349 15614 15355 15631
rect 15326 15611 15355 15614
rect 18315 15610 18318 15636
rect 18344 15610 18347 15636
rect 20064 15631 20093 15634
rect 20064 15630 20070 15631
rect 19198 15616 20070 15630
rect 10243 15563 10272 15566
rect 10243 15546 10249 15563
rect 10266 15562 10272 15563
rect 10449 15562 10452 15568
rect 10266 15548 10452 15562
rect 10266 15546 10272 15548
rect 10243 15543 10272 15546
rect 10449 15542 10452 15548
rect 10478 15542 10481 15568
rect 13509 15563 13538 15566
rect 13509 15546 13515 15563
rect 13532 15562 13538 15563
rect 13669 15562 13672 15568
rect 13532 15548 13672 15562
rect 13532 15546 13538 15548
rect 13509 15543 13538 15546
rect 13669 15542 13672 15548
rect 13698 15542 13701 15568
rect 16245 15542 16248 15568
rect 16274 15562 16277 15568
rect 16361 15563 16390 15566
rect 16361 15562 16367 15563
rect 16274 15548 16367 15562
rect 16274 15542 16277 15548
rect 16361 15546 16367 15548
rect 16384 15546 16390 15563
rect 16361 15543 16390 15546
rect 18315 15542 18318 15568
rect 18344 15562 18347 15568
rect 19198 15562 19212 15616
rect 20064 15614 20070 15616
rect 20087 15614 20093 15631
rect 20064 15611 20093 15614
rect 18344 15548 19212 15562
rect 19351 15563 19380 15566
rect 18344 15542 18347 15548
rect 19351 15546 19357 15563
rect 19374 15562 19380 15563
rect 19971 15562 19974 15568
rect 19374 15548 19974 15562
rect 19374 15546 19380 15548
rect 19351 15543 19380 15546
rect 19971 15542 19974 15548
rect 20000 15542 20003 15568
rect 20072 15562 20086 15611
rect 21029 15610 21032 15636
rect 21058 15610 21061 15636
rect 21397 15610 21400 15636
rect 21426 15630 21429 15636
rect 21797 15630 21811 15645
rect 21903 15644 21906 15645
rect 21932 15644 21935 15670
rect 25353 15644 25356 15670
rect 25382 15644 25385 15670
rect 25523 15668 25537 15684
rect 25565 15682 25571 15699
rect 25565 15679 25586 15682
rect 25583 15678 25586 15679
rect 25612 15678 25615 15704
rect 27299 15670 27328 15671
rect 25515 15665 25544 15668
rect 25515 15648 25521 15665
rect 25538 15664 25544 15665
rect 26043 15664 26046 15670
rect 25538 15650 26046 15664
rect 25538 15648 25544 15650
rect 25515 15645 25544 15648
rect 26043 15644 26046 15650
rect 26072 15644 26075 15670
rect 26917 15644 26920 15670
rect 26946 15664 26949 15670
rect 27101 15664 27104 15670
rect 26946 15650 27104 15664
rect 26946 15644 26949 15650
rect 27101 15644 27104 15650
rect 27130 15664 27133 15670
rect 27148 15665 27177 15668
rect 27148 15664 27154 15665
rect 27130 15650 27154 15664
rect 27130 15644 27133 15650
rect 27148 15648 27154 15650
rect 27171 15648 27177 15665
rect 27148 15645 27177 15648
rect 27193 15644 27196 15670
rect 27222 15668 27225 15670
rect 27222 15665 27234 15668
rect 27228 15648 27234 15665
rect 27222 15645 27234 15648
rect 27222 15644 27225 15645
rect 27285 15644 27288 15670
rect 27314 15668 27328 15670
rect 27322 15651 27328 15668
rect 27314 15648 27328 15651
rect 27314 15644 27317 15648
rect 27346 15644 27349 15670
rect 27375 15644 27378 15670
rect 27409 15665 27438 15668
rect 27409 15648 27415 15665
rect 27432 15664 27438 15665
rect 27460 15665 27489 15668
rect 27432 15648 27446 15664
rect 27409 15645 27446 15648
rect 27460 15648 27466 15665
rect 27483 15664 27489 15665
rect 27561 15664 27564 15670
rect 27483 15650 27564 15664
rect 27483 15648 27489 15650
rect 27460 15645 27489 15648
rect 21426 15616 21811 15630
rect 27432 15630 27446 15645
rect 27561 15644 27564 15650
rect 27590 15644 27593 15670
rect 27745 15630 27748 15636
rect 27432 15616 27748 15630
rect 21426 15610 21429 15616
rect 27745 15610 27748 15616
rect 27774 15610 27777 15636
rect 26503 15576 26506 15602
rect 26532 15596 26535 15602
rect 28113 15596 28116 15602
rect 26532 15582 28116 15596
rect 26532 15576 26535 15582
rect 28113 15576 28116 15582
rect 28142 15576 28145 15602
rect 20247 15562 20250 15568
rect 20072 15548 20250 15562
rect 20247 15542 20250 15548
rect 20276 15542 20279 15568
rect 20293 15542 20296 15568
rect 20322 15562 20325 15568
rect 20385 15562 20388 15568
rect 20322 15548 20388 15562
rect 20322 15542 20325 15548
rect 20385 15542 20388 15548
rect 20414 15542 20417 15568
rect 21582 15563 21611 15566
rect 21582 15546 21588 15563
rect 21605 15562 21611 15563
rect 22823 15562 22826 15568
rect 21605 15548 22826 15562
rect 21605 15546 21611 15548
rect 21582 15543 21611 15546
rect 22823 15542 22826 15548
rect 22852 15542 22855 15568
rect 25997 15542 26000 15568
rect 26026 15562 26029 15568
rect 26319 15562 26322 15568
rect 26026 15548 26322 15562
rect 26026 15542 26029 15548
rect 26319 15542 26322 15548
rect 26348 15542 26351 15568
rect 27101 15542 27104 15568
rect 27130 15562 27133 15568
rect 27331 15562 27334 15568
rect 27130 15548 27334 15562
rect 27130 15542 27133 15548
rect 27331 15542 27334 15548
rect 27360 15542 27363 15568
rect 3036 15480 29992 15528
rect 5711 15460 5714 15466
rect 5582 15446 5714 15460
rect 5582 15396 5596 15446
rect 5711 15440 5714 15446
rect 5740 15440 5743 15466
rect 15923 15440 15926 15466
rect 15952 15460 15955 15466
rect 16429 15460 16432 15466
rect 15952 15446 16432 15460
rect 15952 15440 15955 15446
rect 16429 15440 16432 15446
rect 16458 15440 16461 15466
rect 16935 15440 16938 15466
rect 16964 15460 16967 15466
rect 17971 15461 18000 15464
rect 16964 15446 17924 15460
rect 16964 15440 16967 15446
rect 15932 15426 15946 15440
rect 15886 15412 15946 15426
rect 5574 15393 5603 15396
rect 5574 15376 5580 15393
rect 5597 15376 5603 15393
rect 5574 15373 5603 15376
rect 10771 15372 10774 15398
rect 10800 15392 10803 15398
rect 10864 15393 10893 15396
rect 10864 15392 10870 15393
rect 10800 15378 10870 15392
rect 10800 15372 10803 15378
rect 10864 15376 10870 15378
rect 10887 15376 10893 15393
rect 10864 15373 10893 15376
rect 5619 15338 5622 15364
rect 5648 15358 5651 15364
rect 5735 15359 5764 15362
rect 5735 15358 5741 15359
rect 5648 15344 5741 15358
rect 5648 15338 5651 15344
rect 5735 15342 5741 15344
rect 5758 15358 5764 15359
rect 5987 15358 5990 15364
rect 5758 15344 5990 15358
rect 5758 15342 5764 15344
rect 5735 15339 5764 15342
rect 5987 15338 5990 15344
rect 6016 15338 6019 15364
rect 7275 15338 7278 15364
rect 7304 15358 7307 15364
rect 7413 15358 7416 15364
rect 7304 15344 7416 15358
rect 7304 15338 7307 15344
rect 7413 15338 7416 15344
rect 7442 15358 7445 15364
rect 7828 15359 7857 15362
rect 7828 15358 7834 15359
rect 7442 15344 7834 15358
rect 7442 15338 7445 15344
rect 7828 15342 7834 15344
rect 7851 15342 7857 15359
rect 7828 15339 7857 15342
rect 7989 15359 8018 15362
rect 7989 15342 7995 15359
rect 8012 15358 8018 15359
rect 8103 15358 8106 15364
rect 8012 15344 8106 15358
rect 8012 15342 8018 15344
rect 7989 15339 8018 15342
rect 5785 15325 5814 15328
rect 5785 15308 5791 15325
rect 5808 15324 5814 15325
rect 5849 15324 5852 15330
rect 5808 15310 5852 15324
rect 5808 15308 5814 15310
rect 5785 15305 5814 15308
rect 5849 15304 5852 15310
rect 5878 15304 5881 15330
rect 6999 15304 7002 15330
rect 7028 15324 7031 15330
rect 7091 15324 7094 15330
rect 7028 15310 7094 15324
rect 7028 15304 7031 15310
rect 7091 15304 7094 15310
rect 7120 15304 7123 15330
rect 7781 15304 7784 15330
rect 7810 15324 7813 15330
rect 7997 15324 8011 15339
rect 8103 15338 8106 15344
rect 8132 15338 8135 15364
rect 8425 15358 8428 15364
rect 8158 15344 8428 15358
rect 7810 15310 8011 15324
rect 8039 15325 8068 15328
rect 7810 15304 7813 15310
rect 8039 15308 8045 15325
rect 8062 15324 8068 15325
rect 8158 15324 8172 15344
rect 8425 15338 8428 15344
rect 8454 15338 8457 15364
rect 10909 15338 10912 15364
rect 10938 15358 10941 15364
rect 11019 15359 11048 15362
rect 11019 15358 11025 15359
rect 10938 15344 11025 15358
rect 10938 15338 10941 15344
rect 11019 15342 11025 15344
rect 11042 15358 11048 15359
rect 11139 15358 11142 15364
rect 11042 15344 11142 15358
rect 11042 15342 11048 15344
rect 11019 15339 11048 15342
rect 11139 15338 11142 15344
rect 11168 15338 11171 15364
rect 13255 15338 13258 15364
rect 13284 15358 13287 15364
rect 13807 15358 13810 15364
rect 13284 15344 13810 15358
rect 13284 15338 13287 15344
rect 13807 15338 13810 15344
rect 13836 15338 13839 15364
rect 13945 15338 13948 15364
rect 13974 15362 13977 15364
rect 15886 15362 15900 15412
rect 15924 15393 15953 15396
rect 15924 15376 15930 15393
rect 15947 15392 15953 15393
rect 16061 15392 16064 15398
rect 15947 15378 16064 15392
rect 15947 15376 15953 15378
rect 15924 15373 15953 15376
rect 16061 15372 16064 15378
rect 16090 15372 16093 15398
rect 16153 15372 16156 15398
rect 16182 15392 16185 15398
rect 16246 15393 16275 15396
rect 16246 15392 16252 15393
rect 16182 15378 16252 15392
rect 16182 15372 16185 15378
rect 16246 15376 16252 15378
rect 16269 15376 16275 15393
rect 17910 15392 17924 15446
rect 17971 15444 17977 15461
rect 17994 15460 18000 15461
rect 18913 15460 18916 15466
rect 17994 15446 18916 15460
rect 17994 15444 18000 15446
rect 17971 15441 18000 15444
rect 18913 15440 18916 15446
rect 18942 15440 18945 15466
rect 20063 15440 20066 15466
rect 20092 15460 20095 15466
rect 22639 15460 22642 15466
rect 20092 15446 22642 15460
rect 20092 15440 20095 15446
rect 22639 15440 22642 15446
rect 22668 15460 22671 15466
rect 25285 15461 25314 15464
rect 22668 15446 25238 15460
rect 22668 15440 22671 15446
rect 20201 15406 20204 15432
rect 20230 15426 20233 15432
rect 25224 15426 25238 15446
rect 25285 15444 25291 15461
rect 25308 15460 25314 15461
rect 25675 15460 25678 15466
rect 25308 15446 25678 15460
rect 25308 15444 25314 15446
rect 25285 15441 25314 15444
rect 25675 15440 25678 15446
rect 25704 15440 25707 15466
rect 27745 15440 27748 15466
rect 27774 15464 27777 15466
rect 27774 15461 27798 15464
rect 27774 15444 27775 15461
rect 27792 15444 27798 15461
rect 27774 15441 27798 15444
rect 27774 15440 27777 15441
rect 25721 15426 25724 15432
rect 20230 15412 20408 15426
rect 25224 15412 25724 15426
rect 20230 15406 20233 15412
rect 18315 15392 18318 15398
rect 17910 15378 18318 15392
rect 16246 15373 16275 15376
rect 18315 15372 18318 15378
rect 18344 15392 18347 15398
rect 18454 15393 18483 15396
rect 18454 15392 18460 15393
rect 18344 15378 18460 15392
rect 18344 15372 18347 15378
rect 18454 15376 18460 15378
rect 18477 15376 18483 15393
rect 18454 15373 18483 15376
rect 20064 15393 20093 15396
rect 20064 15376 20070 15393
rect 20087 15392 20093 15393
rect 20087 15378 20362 15392
rect 20087 15376 20093 15378
rect 20064 15373 20093 15376
rect 13974 15359 13992 15362
rect 13986 15342 13992 15359
rect 13974 15339 13992 15342
rect 15878 15359 15907 15362
rect 15878 15342 15884 15359
rect 15901 15342 15907 15359
rect 15878 15339 15907 15342
rect 13974 15338 13977 15339
rect 15969 15338 15972 15364
rect 15998 15362 16001 15364
rect 15998 15358 16002 15362
rect 15998 15344 16020 15358
rect 15998 15339 16002 15344
rect 15998 15338 16001 15339
rect 16107 15338 16110 15364
rect 16136 15358 16139 15364
rect 16433 15359 16462 15362
rect 16433 15358 16439 15359
rect 16136 15344 16439 15358
rect 16136 15338 16139 15344
rect 16433 15342 16439 15344
rect 16456 15358 16462 15359
rect 16889 15358 16892 15364
rect 16456 15344 16892 15358
rect 16456 15342 16462 15344
rect 16433 15339 16462 15342
rect 16889 15338 16892 15344
rect 16918 15338 16921 15364
rect 16935 15338 16938 15364
rect 16964 15338 16967 15364
rect 18615 15359 18644 15362
rect 18615 15342 18621 15359
rect 18638 15358 18644 15359
rect 18729 15358 18732 15364
rect 18638 15344 18732 15358
rect 18638 15342 18644 15344
rect 18615 15339 18644 15342
rect 18729 15338 18732 15344
rect 18758 15338 18761 15364
rect 18867 15358 18870 15364
rect 18784 15344 18870 15358
rect 11093 15328 11096 15330
rect 8062 15310 8172 15324
rect 11075 15325 11096 15328
rect 8062 15308 8068 15310
rect 8039 15305 8068 15308
rect 11075 15308 11081 15325
rect 11075 15305 11096 15308
rect 11093 15304 11096 15305
rect 11122 15304 11125 15330
rect 14037 15328 14040 15330
rect 14019 15325 14040 15328
rect 14019 15308 14025 15325
rect 14019 15305 14040 15308
rect 14037 15304 14040 15305
rect 14066 15304 14069 15330
rect 15785 15304 15788 15330
rect 15814 15304 15817 15330
rect 15924 15325 15953 15328
rect 15924 15308 15930 15325
rect 15947 15324 15953 15325
rect 16199 15324 16202 15330
rect 15947 15310 16202 15324
rect 15947 15308 15953 15310
rect 15924 15305 15953 15308
rect 16199 15304 16202 15310
rect 16228 15304 16231 15330
rect 16245 15304 16248 15330
rect 16274 15304 16277 15330
rect 16337 15304 16340 15330
rect 16366 15304 16369 15330
rect 16383 15304 16386 15330
rect 16412 15304 16415 15330
rect 16567 15304 16570 15330
rect 16596 15324 16599 15330
rect 17165 15328 17168 15330
rect 17096 15325 17125 15328
rect 17096 15324 17102 15325
rect 16596 15310 17102 15324
rect 16596 15304 16599 15310
rect 17096 15308 17102 15310
rect 17119 15308 17125 15325
rect 17096 15305 17125 15308
rect 17147 15325 17168 15328
rect 17147 15308 17153 15325
rect 17147 15305 17168 15308
rect 17165 15304 17168 15305
rect 17194 15304 17197 15330
rect 18683 15328 18686 15330
rect 18665 15325 18686 15328
rect 18665 15308 18671 15325
rect 18712 15324 18715 15330
rect 18784 15324 18798 15344
rect 18867 15338 18870 15344
rect 18896 15338 18899 15364
rect 19489 15359 19518 15362
rect 19489 15342 19495 15359
rect 19512 15358 19518 15359
rect 20110 15359 20139 15362
rect 20110 15358 20116 15359
rect 19512 15344 20116 15358
rect 19512 15342 19518 15344
rect 19489 15339 19518 15342
rect 20110 15342 20116 15344
rect 20133 15342 20139 15359
rect 20110 15339 20139 15342
rect 20159 15359 20188 15362
rect 20159 15342 20165 15359
rect 20182 15342 20188 15359
rect 20159 15339 20188 15342
rect 18712 15310 18798 15324
rect 18665 15305 18686 15308
rect 18683 15304 18686 15305
rect 18712 15304 18715 15310
rect 19971 15304 19974 15330
rect 20000 15304 20003 15330
rect 20063 15304 20066 15330
rect 20092 15304 20095 15330
rect 20164 15324 20178 15339
rect 20201 15324 20204 15330
rect 20164 15310 20204 15324
rect 20201 15304 20204 15310
rect 20230 15304 20233 15330
rect 20348 15324 20362 15378
rect 20394 15358 20408 15412
rect 25721 15406 25724 15412
rect 25750 15406 25753 15432
rect 22823 15372 22826 15398
rect 22852 15372 22855 15398
rect 24157 15372 24160 15398
rect 24186 15392 24189 15398
rect 24250 15393 24279 15396
rect 24250 15392 24256 15393
rect 24186 15378 24256 15392
rect 24186 15372 24189 15378
rect 24250 15376 24256 15378
rect 24273 15376 24279 15393
rect 24250 15373 24279 15376
rect 26733 15372 26736 15398
rect 26762 15372 26765 15398
rect 20937 15358 20940 15364
rect 20394 15344 20940 15358
rect 20937 15338 20940 15344
rect 20966 15338 20969 15364
rect 22732 15359 22761 15362
rect 22732 15342 22738 15359
rect 22755 15358 22761 15359
rect 22869 15358 22872 15364
rect 22755 15344 22872 15358
rect 22755 15342 22761 15344
rect 22732 15339 22761 15342
rect 22869 15338 22872 15344
rect 22898 15338 22901 15364
rect 22915 15338 22918 15364
rect 22944 15338 22947 15364
rect 24387 15338 24390 15364
rect 24416 15362 24419 15364
rect 24416 15359 24434 15362
rect 24428 15342 24434 15359
rect 24416 15339 24434 15342
rect 24416 15338 24419 15339
rect 26779 15338 26782 15364
rect 26808 15358 26811 15364
rect 26889 15359 26918 15362
rect 26889 15358 26895 15359
rect 26808 15344 26895 15358
rect 26808 15338 26811 15344
rect 26889 15342 26895 15344
rect 26912 15342 26918 15359
rect 26889 15339 26918 15342
rect 22778 15325 22807 15328
rect 22778 15324 22784 15325
rect 20348 15310 22784 15324
rect 22778 15308 22784 15310
rect 22801 15308 22807 15325
rect 22778 15305 22807 15308
rect 22961 15304 22964 15330
rect 22990 15324 22993 15330
rect 26963 15328 26966 15330
rect 24449 15325 24478 15328
rect 24449 15324 24455 15325
rect 22990 15310 24455 15324
rect 22990 15304 22993 15310
rect 24449 15308 24455 15310
rect 24472 15308 24478 15325
rect 24449 15305 24478 15308
rect 26945 15325 26966 15328
rect 26945 15308 26951 15325
rect 26945 15305 26966 15308
rect 26963 15304 26966 15305
rect 26992 15304 26995 15330
rect 6609 15291 6638 15294
rect 6609 15274 6615 15291
rect 6632 15290 6638 15291
rect 6769 15290 6772 15296
rect 6632 15276 6772 15290
rect 6632 15274 6638 15276
rect 6609 15271 6638 15274
rect 6769 15270 6772 15276
rect 6798 15270 6801 15296
rect 8863 15291 8892 15294
rect 8863 15274 8869 15291
rect 8886 15290 8892 15291
rect 9069 15290 9072 15296
rect 8886 15276 9072 15290
rect 8886 15274 8892 15276
rect 8863 15271 8892 15274
rect 9069 15270 9072 15276
rect 9098 15270 9101 15296
rect 11899 15291 11928 15294
rect 11899 15274 11905 15291
rect 11922 15290 11928 15291
rect 11967 15290 11970 15296
rect 11922 15276 11970 15290
rect 11922 15274 11928 15276
rect 11899 15271 11928 15274
rect 11967 15270 11970 15276
rect 11996 15270 11999 15296
rect 14819 15270 14822 15296
rect 14848 15294 14851 15296
rect 14848 15291 14872 15294
rect 14848 15274 14849 15291
rect 14866 15274 14872 15291
rect 14848 15271 14872 15274
rect 14848 15270 14851 15271
rect 22869 15270 22872 15296
rect 22898 15270 22901 15296
rect 3036 15208 29992 15256
rect 5941 15168 5944 15194
rect 5970 15188 5973 15194
rect 6448 15189 6477 15192
rect 6448 15188 6454 15189
rect 5970 15174 6454 15188
rect 5970 15168 5973 15174
rect 6448 15172 6454 15174
rect 6471 15172 6477 15189
rect 7137 15188 7140 15194
rect 6448 15169 6477 15172
rect 7008 15174 7140 15188
rect 3779 15158 3782 15160
rect 3761 15155 3782 15158
rect 3761 15138 3767 15155
rect 3761 15135 3782 15138
rect 3779 15134 3782 15135
rect 3808 15134 3811 15160
rect 4930 15155 4959 15158
rect 4930 15138 4936 15155
rect 4953 15154 4959 15155
rect 5159 15154 5162 15160
rect 4953 15140 5162 15154
rect 4953 15138 4959 15140
rect 4930 15135 4959 15138
rect 5159 15134 5162 15140
rect 5188 15134 5191 15160
rect 6861 15134 6864 15160
rect 6890 15134 6893 15160
rect 7008 15154 7022 15174
rect 7137 15168 7140 15174
rect 7166 15168 7169 15194
rect 8977 15188 8980 15194
rect 8940 15174 8980 15188
rect 6962 15140 7022 15154
rect 3411 15100 3414 15126
rect 3440 15120 3443 15126
rect 3705 15121 3734 15124
rect 3705 15120 3711 15121
rect 3440 15106 3711 15120
rect 3440 15100 3443 15106
rect 3705 15104 3711 15106
rect 3728 15104 3734 15121
rect 3705 15101 3734 15104
rect 4837 15100 4840 15126
rect 4866 15100 4869 15126
rect 4975 15100 4978 15126
rect 5004 15100 5007 15126
rect 5022 15121 5051 15124
rect 5022 15104 5028 15121
rect 5045 15120 5051 15121
rect 5067 15120 5070 15126
rect 5045 15106 5070 15120
rect 5045 15104 5051 15106
rect 5022 15101 5051 15104
rect 5067 15100 5070 15106
rect 5096 15100 5099 15126
rect 6356 15121 6385 15124
rect 6356 15104 6362 15121
rect 6379 15104 6385 15121
rect 6356 15101 6385 15104
rect 6402 15121 6431 15124
rect 6402 15104 6408 15121
rect 6425 15120 6431 15121
rect 6447 15120 6450 15126
rect 6425 15106 6450 15120
rect 6425 15104 6431 15106
rect 6402 15101 6431 15104
rect 3457 15066 3460 15092
rect 3486 15086 3489 15092
rect 3550 15087 3579 15090
rect 3550 15086 3556 15087
rect 3486 15072 3556 15086
rect 3486 15066 3489 15072
rect 3550 15070 3556 15072
rect 3573 15070 3579 15087
rect 6364 15086 6378 15101
rect 6447 15100 6450 15106
rect 6476 15100 6479 15126
rect 6540 15121 6569 15124
rect 6540 15104 6546 15121
rect 6563 15120 6569 15121
rect 6631 15120 6634 15126
rect 6563 15106 6634 15120
rect 6563 15104 6569 15106
rect 6540 15101 6569 15104
rect 6631 15100 6634 15106
rect 6660 15100 6663 15126
rect 6769 15100 6772 15126
rect 6798 15100 6801 15126
rect 6907 15100 6910 15126
rect 6936 15100 6939 15126
rect 6962 15124 6976 15140
rect 7045 15134 7048 15160
rect 7074 15154 7077 15160
rect 7436 15155 7465 15158
rect 7074 15140 7390 15154
rect 7074 15134 7077 15140
rect 6954 15121 6983 15124
rect 6954 15104 6960 15121
rect 6977 15104 6983 15121
rect 7321 15120 7324 15126
rect 6954 15101 6983 15104
rect 7008 15106 7324 15120
rect 7008 15086 7022 15106
rect 7321 15100 7324 15106
rect 7350 15100 7353 15126
rect 7376 15120 7390 15140
rect 7436 15138 7442 15155
rect 7459 15154 7465 15155
rect 8940 15154 8954 15174
rect 8977 15168 8980 15174
rect 9006 15168 9009 15194
rect 9069 15188 9072 15194
rect 9063 15168 9072 15188
rect 9098 15168 9101 15194
rect 10541 15168 10544 15194
rect 10570 15188 10573 15194
rect 10570 15174 11927 15188
rect 10570 15168 10573 15174
rect 7459 15140 7574 15154
rect 7459 15138 7465 15140
rect 7436 15135 7465 15138
rect 7475 15121 7504 15124
rect 7475 15120 7481 15121
rect 7376 15106 7481 15120
rect 7475 15104 7481 15106
rect 7498 15104 7504 15121
rect 7560 15120 7574 15140
rect 8802 15140 8954 15154
rect 7827 15120 7830 15126
rect 7560 15106 7830 15120
rect 7475 15101 7504 15104
rect 7827 15100 7830 15106
rect 7856 15100 7859 15126
rect 8802 15124 8816 15140
rect 9063 15135 9077 15168
rect 10265 15158 10268 15160
rect 10243 15155 10268 15158
rect 10243 15154 10249 15155
rect 9262 15140 10249 15154
rect 9055 15132 9084 15135
rect 8794 15121 8823 15124
rect 8794 15104 8800 15121
rect 8817 15104 8823 15121
rect 8794 15101 8823 15104
rect 8839 15100 8842 15126
rect 8868 15124 8871 15126
rect 8868 15121 8880 15124
rect 8874 15104 8880 15121
rect 8945 15121 8974 15124
rect 8945 15120 8951 15121
rect 8868 15101 8880 15104
rect 8940 15104 8951 15120
rect 8968 15104 8974 15121
rect 8940 15101 8974 15104
rect 9007 15121 9036 15124
rect 9007 15104 9013 15121
rect 9030 15104 9036 15121
rect 9055 15115 9061 15132
rect 9078 15115 9084 15132
rect 9055 15112 9084 15115
rect 9106 15121 9135 15124
rect 9007 15101 9036 15104
rect 9106 15104 9112 15121
rect 9129 15120 9135 15121
rect 9207 15120 9210 15126
rect 9129 15106 9210 15120
rect 9129 15104 9135 15106
rect 9106 15101 9135 15104
rect 8868 15100 8871 15101
rect 6364 15072 7022 15086
rect 3550 15067 3579 15070
rect 7275 15066 7278 15092
rect 7304 15066 7307 15092
rect 8311 15087 8340 15090
rect 8311 15070 8317 15087
rect 8334 15086 8340 15087
rect 8940 15086 8954 15101
rect 8334 15072 8954 15086
rect 9015 15086 9029 15101
rect 9207 15100 9210 15106
rect 9236 15100 9239 15126
rect 9161 15086 9164 15092
rect 9015 15072 9164 15086
rect 8334 15070 8340 15072
rect 8311 15067 8340 15070
rect 9161 15066 9164 15072
rect 9190 15066 9193 15092
rect 4699 15032 4702 15058
rect 4728 15052 4731 15058
rect 5021 15052 5024 15058
rect 4728 15038 5024 15052
rect 4728 15032 4731 15038
rect 5021 15032 5024 15038
rect 5050 15032 5053 15058
rect 8885 15032 8888 15058
rect 8914 15052 8917 15058
rect 9262 15052 9276 15140
rect 10243 15138 10249 15140
rect 10266 15138 10268 15155
rect 10243 15135 10268 15138
rect 10265 15134 10268 15135
rect 10294 15134 10297 15160
rect 11071 15155 11100 15158
rect 11071 15138 11077 15155
rect 11094 15154 11100 15155
rect 11094 15140 11760 15154
rect 11094 15138 11100 15140
rect 11071 15135 11100 15138
rect 10197 15121 10226 15124
rect 10197 15104 10203 15121
rect 10220 15120 10226 15121
rect 10909 15120 10912 15126
rect 10220 15106 10912 15120
rect 10220 15104 10226 15106
rect 10197 15101 10226 15104
rect 10909 15100 10912 15106
rect 10938 15100 10941 15126
rect 11746 15124 11760 15140
rect 11692 15121 11721 15124
rect 11692 15104 11698 15121
rect 11715 15104 11721 15121
rect 11746 15121 11778 15124
rect 11746 15106 11755 15121
rect 11692 15101 11721 15104
rect 11749 15104 11755 15106
rect 11772 15104 11778 15121
rect 11749 15101 11778 15104
rect 10036 15087 10065 15090
rect 10036 15086 10042 15087
rect 8914 15038 9276 15052
rect 9653 15072 10042 15086
rect 8914 15032 8917 15038
rect 4585 15019 4614 15022
rect 4585 15002 4591 15019
rect 4608 15018 4614 15019
rect 4791 15018 4794 15024
rect 4608 15004 4794 15018
rect 4608 15002 4614 15004
rect 4585 14999 4614 15002
rect 4791 14998 4794 15004
rect 4820 14998 4823 15024
rect 5113 14998 5116 15024
rect 5142 14998 5145 15024
rect 6401 14998 6404 15024
rect 6430 14998 6433 15024
rect 7046 15019 7075 15022
rect 7046 15002 7052 15019
rect 7069 15018 7075 15019
rect 7413 15018 7416 15024
rect 7069 15004 7416 15018
rect 7069 15002 7075 15004
rect 7046 14999 7075 15002
rect 7413 14998 7416 15004
rect 7442 14998 7445 15024
rect 7459 14998 7462 15024
rect 7488 15018 7491 15024
rect 8794 15019 8823 15022
rect 8794 15018 8800 15019
rect 7488 15004 8800 15018
rect 7488 14998 7491 15004
rect 8794 15002 8800 15004
rect 8817 15002 8823 15019
rect 8794 14999 8823 15002
rect 9115 14998 9118 15024
rect 9144 15018 9147 15024
rect 9653 15018 9667 15072
rect 10036 15070 10042 15072
rect 10059 15070 10065 15087
rect 10036 15067 10065 15070
rect 11700 15052 11714 15101
rect 11829 15100 11832 15126
rect 11858 15124 11861 15126
rect 11913 15124 11927 15174
rect 11967 15168 11970 15194
rect 11996 15168 11999 15194
rect 16383 15168 16386 15194
rect 16412 15192 16415 15194
rect 16412 15189 16436 15192
rect 16412 15172 16413 15189
rect 16430 15172 16436 15189
rect 16412 15169 16436 15172
rect 21559 15189 21588 15192
rect 21559 15172 21565 15189
rect 21582 15188 21588 15189
rect 21719 15188 21722 15194
rect 21582 15174 21722 15188
rect 21582 15172 21588 15174
rect 21559 15169 21588 15172
rect 16412 15168 16415 15169
rect 21719 15168 21722 15174
rect 21748 15168 21751 15194
rect 11976 15124 11990 15168
rect 12841 15134 12844 15160
rect 12870 15154 12873 15160
rect 13025 15158 13028 15160
rect 12956 15155 12985 15158
rect 12956 15154 12962 15155
rect 12870 15140 12962 15154
rect 12870 15134 12873 15140
rect 12956 15138 12962 15140
rect 12979 15138 12985 15155
rect 12956 15135 12985 15138
rect 13007 15155 13028 15158
rect 13007 15138 13013 15155
rect 13007 15135 13028 15138
rect 13025 15134 13028 15135
rect 13054 15134 13057 15160
rect 13831 15155 13860 15158
rect 13831 15138 13837 15155
rect 13854 15154 13860 15155
rect 14819 15154 14822 15160
rect 13854 15140 14612 15154
rect 13854 15138 13860 15140
rect 13831 15135 13860 15138
rect 14598 15127 14612 15140
rect 14736 15140 14822 15154
rect 11858 15121 11872 15124
rect 11866 15104 11872 15121
rect 11858 15101 11872 15104
rect 11905 15121 11934 15124
rect 11905 15104 11911 15121
rect 11928 15104 11934 15121
rect 11905 15101 11934 15104
rect 11953 15121 11990 15124
rect 11953 15104 11959 15121
rect 11976 15106 11990 15121
rect 12004 15124 12033 15127
rect 12004 15107 12010 15124
rect 12027 15120 12033 15124
rect 12059 15120 12062 15126
rect 12027 15107 12062 15120
rect 12004 15106 12062 15107
rect 11976 15104 11982 15106
rect 12004 15104 12033 15106
rect 11953 15101 11982 15104
rect 11858 15100 11861 15101
rect 11913 15086 11927 15101
rect 12059 15100 12062 15106
rect 12088 15120 12091 15126
rect 14452 15121 14481 15124
rect 14452 15120 14458 15121
rect 12088 15106 13738 15120
rect 12088 15100 12091 15106
rect 13724 15092 13738 15106
rect 13770 15106 14458 15120
rect 12105 15086 12108 15092
rect 11913 15072 12108 15086
rect 12105 15066 12108 15072
rect 12134 15066 12137 15092
rect 12381 15066 12384 15092
rect 12410 15086 12413 15092
rect 12796 15087 12825 15090
rect 12796 15086 12802 15087
rect 12410 15072 12802 15086
rect 12410 15066 12413 15072
rect 12796 15070 12802 15072
rect 12819 15070 12825 15087
rect 12796 15067 12825 15070
rect 13715 15066 13718 15092
rect 13744 15066 13747 15092
rect 11033 15038 12082 15052
rect 9144 15004 9667 15018
rect 9144 14998 9147 15004
rect 10173 14998 10176 15024
rect 10202 15018 10205 15024
rect 11033 15018 11047 15038
rect 10202 15004 11047 15018
rect 11692 15019 11721 15022
rect 10202 14998 10205 15004
rect 11692 15002 11698 15019
rect 11715 15018 11721 15019
rect 12013 15018 12016 15024
rect 11715 15004 12016 15018
rect 11715 15002 11721 15004
rect 11692 14999 11721 15002
rect 12013 14998 12016 15004
rect 12042 14998 12045 15024
rect 12068 15018 12082 15038
rect 13393 15018 13396 15024
rect 12068 15004 13396 15018
rect 13393 14998 13396 15004
rect 13422 15018 13425 15024
rect 13770 15018 13784 15106
rect 14452 15104 14458 15106
rect 14475 15104 14481 15121
rect 14452 15101 14481 15104
rect 14497 15100 14500 15126
rect 14526 15124 14529 15126
rect 14598 15124 14632 15127
rect 14526 15121 14538 15124
rect 14532 15104 14538 15121
rect 14598 15107 14609 15124
rect 14626 15107 14632 15124
rect 14736 15119 14750 15140
rect 14819 15134 14822 15140
rect 14848 15134 14851 15160
rect 15279 15134 15282 15160
rect 15308 15154 15311 15160
rect 15601 15158 15604 15160
rect 15583 15155 15604 15158
rect 15583 15154 15589 15155
rect 15308 15140 15589 15154
rect 15308 15134 15311 15140
rect 15583 15138 15589 15140
rect 15583 15135 15604 15138
rect 15601 15134 15604 15135
rect 15630 15134 15633 15160
rect 20753 15158 20756 15160
rect 20735 15155 20756 15158
rect 20735 15138 20741 15155
rect 20735 15135 20756 15138
rect 20753 15134 20756 15135
rect 20782 15134 20785 15160
rect 28389 15134 28392 15160
rect 28418 15154 28421 15160
rect 28573 15158 28576 15160
rect 28551 15155 28576 15158
rect 28551 15154 28557 15155
rect 28418 15140 28557 15154
rect 28418 15134 28421 15140
rect 28551 15138 28557 15140
rect 28574 15138 28576 15155
rect 28551 15135 28576 15138
rect 28573 15134 28576 15135
rect 28602 15134 28605 15160
rect 14598 15106 14632 15107
rect 14603 15104 14632 15106
rect 14651 15116 14680 15119
rect 14526 15101 14538 15104
rect 14526 15100 14529 15101
rect 14651 15099 14657 15116
rect 14674 15099 14680 15116
rect 14651 15096 14680 15099
rect 14713 15116 14750 15119
rect 14713 15099 14719 15116
rect 14736 15100 14750 15116
rect 14764 15121 14793 15124
rect 14764 15104 14770 15121
rect 14787 15120 14793 15121
rect 15233 15120 15236 15126
rect 14787 15106 15236 15120
rect 14787 15104 14793 15106
rect 14764 15101 14793 15104
rect 15233 15100 15236 15106
rect 15262 15100 15265 15126
rect 15509 15100 15512 15126
rect 15538 15124 15541 15126
rect 15538 15121 15556 15124
rect 15550 15104 15556 15121
rect 15538 15101 15556 15104
rect 15538 15100 15541 15101
rect 18407 15100 18410 15126
rect 18436 15120 18439 15126
rect 18500 15121 18529 15124
rect 18500 15120 18506 15121
rect 18436 15106 18506 15120
rect 18436 15100 18439 15106
rect 18500 15104 18506 15106
rect 18523 15104 18529 15121
rect 18500 15101 18529 15104
rect 18913 15100 18916 15126
rect 18942 15100 18945 15126
rect 20247 15100 20250 15126
rect 20276 15120 20279 15126
rect 20524 15121 20553 15124
rect 20524 15120 20530 15121
rect 20276 15106 20530 15120
rect 20276 15100 20279 15106
rect 20524 15104 20530 15106
rect 20547 15120 20553 15121
rect 20569 15120 20572 15126
rect 20547 15106 20572 15120
rect 20547 15104 20553 15106
rect 20524 15101 20553 15104
rect 20569 15100 20572 15106
rect 20598 15100 20601 15126
rect 20685 15121 20714 15124
rect 20685 15104 20691 15121
rect 20708 15120 20714 15121
rect 20799 15120 20802 15126
rect 20708 15106 20802 15120
rect 20708 15104 20714 15106
rect 20685 15101 20714 15104
rect 20799 15100 20802 15106
rect 20828 15100 20831 15126
rect 28297 15100 28300 15126
rect 28326 15120 28329 15126
rect 28344 15121 28373 15124
rect 28344 15120 28350 15121
rect 28326 15106 28350 15120
rect 28326 15100 28329 15106
rect 28344 15104 28350 15106
rect 28367 15104 28373 15121
rect 28499 15121 28528 15124
rect 28499 15120 28505 15121
rect 28344 15101 28373 15104
rect 28398 15106 28505 15120
rect 14736 15099 14742 15100
rect 14713 15096 14742 15099
rect 14267 15066 14270 15092
rect 14296 15086 14299 15092
rect 14296 15072 14497 15086
rect 14296 15066 14299 15072
rect 14483 15052 14497 15072
rect 14659 15052 14673 15096
rect 15187 15066 15190 15092
rect 15216 15086 15219 15092
rect 15372 15087 15401 15090
rect 15372 15086 15378 15087
rect 15216 15072 15378 15086
rect 15216 15066 15219 15072
rect 15372 15070 15378 15072
rect 15395 15070 15401 15087
rect 15372 15067 15401 15070
rect 18730 15087 18759 15090
rect 18730 15070 18736 15087
rect 18753 15070 18759 15087
rect 28398 15086 28412 15106
rect 28499 15104 28505 15106
rect 28522 15104 28528 15121
rect 28499 15101 28528 15104
rect 18730 15067 18759 15070
rect 28306 15072 28412 15086
rect 14483 15038 14673 15052
rect 13422 15004 13784 15018
rect 14452 15019 14481 15022
rect 13422 14998 13425 15004
rect 14452 15002 14458 15019
rect 14475 15018 14481 15019
rect 16015 15018 16018 15024
rect 14475 15004 16018 15018
rect 14475 15002 14481 15004
rect 14452 14999 14481 15002
rect 16015 14998 16018 15004
rect 16044 14998 16047 15024
rect 18738 15018 18752 15067
rect 28306 15058 28320 15072
rect 21498 15038 25537 15052
rect 21498 15018 21512 15038
rect 18738 15004 21512 15018
rect 25523 15018 25537 15038
rect 28297 15032 28300 15058
rect 28326 15032 28329 15058
rect 31747 15052 31750 15058
rect 29180 15038 31750 15052
rect 29180 15018 29194 15038
rect 31747 15032 31750 15038
rect 31776 15032 31779 15058
rect 25523 15004 29194 15018
rect 29379 15019 29408 15022
rect 29379 15002 29385 15019
rect 29402 15018 29408 15019
rect 29447 15018 29450 15024
rect 29402 15004 29450 15018
rect 29402 15002 29408 15004
rect 29379 14999 29408 15002
rect 29447 14998 29450 15004
rect 29476 14998 29479 15024
rect 3036 14936 29992 14984
rect 3319 14916 3322 14922
rect 3144 14902 3322 14916
rect 3144 14852 3158 14902
rect 3319 14896 3322 14902
rect 3348 14916 3351 14922
rect 3457 14916 3460 14922
rect 3348 14902 3460 14916
rect 3348 14896 3351 14902
rect 3457 14896 3460 14902
rect 3486 14896 3489 14922
rect 4171 14917 4200 14920
rect 4171 14900 4177 14917
rect 4194 14916 4200 14917
rect 4837 14916 4840 14922
rect 4194 14902 4840 14916
rect 4194 14900 4200 14902
rect 4171 14897 4200 14900
rect 4837 14896 4840 14902
rect 4866 14896 4869 14922
rect 6447 14896 6450 14922
rect 6476 14916 6479 14922
rect 7414 14917 7443 14920
rect 7414 14916 7420 14917
rect 6476 14902 7420 14916
rect 6476 14896 6479 14902
rect 7414 14900 7420 14902
rect 7437 14900 7443 14917
rect 7414 14897 7443 14900
rect 9207 14896 9210 14922
rect 9236 14916 9239 14922
rect 12059 14916 12062 14922
rect 9236 14902 12062 14916
rect 9236 14896 9239 14902
rect 10449 14882 10452 14888
rect 10443 14862 10452 14882
rect 10478 14862 10481 14888
rect 3136 14849 3165 14852
rect 3136 14832 3142 14849
rect 3159 14832 3165 14849
rect 5113 14848 5116 14854
rect 3136 14829 3165 14832
rect 4754 14834 5116 14848
rect 3181 14794 3184 14820
rect 3210 14814 3213 14820
rect 4754 14818 4768 14834
rect 5113 14828 5116 14834
rect 5142 14828 5145 14854
rect 6931 14849 6960 14852
rect 6931 14832 6937 14849
rect 6954 14848 6960 14849
rect 6954 14834 7620 14848
rect 6954 14832 6960 14834
rect 6931 14829 6960 14832
rect 4746 14815 4775 14818
rect 3210 14800 3368 14814
rect 3210 14794 3213 14800
rect 3354 14784 3368 14800
rect 4746 14798 4752 14815
rect 4769 14798 4775 14815
rect 4746 14795 4775 14798
rect 4791 14794 4794 14820
rect 4820 14794 4823 14820
rect 4837 14794 4840 14820
rect 4866 14814 4869 14820
rect 4976 14815 5005 14818
rect 4976 14814 4982 14815
rect 4866 14800 4982 14814
rect 4866 14794 4869 14800
rect 4976 14798 4982 14800
rect 4999 14798 5005 14815
rect 4976 14795 5005 14798
rect 5895 14794 5898 14820
rect 5924 14794 5927 14820
rect 6033 14794 6036 14820
rect 6062 14818 6065 14820
rect 6062 14815 6080 14818
rect 6074 14798 6080 14815
rect 6999 14814 7002 14820
rect 6062 14795 6080 14798
rect 6226 14800 7002 14814
rect 6062 14794 6065 14795
rect 3296 14781 3325 14784
rect 3296 14780 3302 14781
rect 3190 14766 3302 14780
rect 3190 14752 3204 14766
rect 3296 14764 3302 14766
rect 3319 14764 3325 14781
rect 3296 14761 3325 14764
rect 3347 14781 3368 14784
rect 3347 14764 3353 14781
rect 3347 14761 3368 14764
rect 3365 14760 3368 14761
rect 3394 14760 3397 14786
rect 4883 14760 4886 14786
rect 4912 14760 4915 14786
rect 4929 14760 4932 14786
rect 4958 14760 4961 14786
rect 6125 14784 6128 14786
rect 6107 14781 6128 14784
rect 6107 14764 6113 14781
rect 6154 14780 6157 14786
rect 6226 14780 6240 14800
rect 6999 14794 7002 14800
rect 7028 14794 7031 14820
rect 7413 14794 7416 14820
rect 7442 14794 7445 14820
rect 7459 14794 7462 14820
rect 7488 14794 7491 14820
rect 7606 14818 7620 14834
rect 10443 14824 10457 14862
rect 10435 14821 10464 14824
rect 7598 14815 7627 14818
rect 7598 14798 7604 14815
rect 7621 14798 7627 14815
rect 7598 14795 7627 14798
rect 7644 14815 7673 14818
rect 7644 14798 7650 14815
rect 7667 14814 7673 14815
rect 7689 14814 7692 14820
rect 7667 14800 7692 14814
rect 7667 14798 7673 14800
rect 7644 14795 7673 14798
rect 7689 14794 7692 14800
rect 7718 14794 7721 14820
rect 8287 14794 8290 14820
rect 8316 14814 8319 14820
rect 8316 14800 8402 14814
rect 8316 14794 8319 14800
rect 6154 14766 6240 14780
rect 7552 14781 7581 14784
rect 6107 14761 6128 14764
rect 6125 14760 6128 14761
rect 6154 14760 6157 14766
rect 7552 14764 7558 14781
rect 7575 14780 7581 14781
rect 8241 14780 8244 14786
rect 7575 14766 8244 14780
rect 7575 14764 7581 14766
rect 7552 14761 7581 14764
rect 8241 14760 8244 14766
rect 8270 14760 8273 14786
rect 8388 14780 8402 14800
rect 8517 14794 8520 14820
rect 8546 14814 8549 14820
rect 8656 14815 8685 14818
rect 8656 14814 8662 14815
rect 8546 14800 8662 14814
rect 8546 14794 8549 14800
rect 8656 14798 8662 14800
rect 8679 14798 8685 14815
rect 8656 14795 8685 14798
rect 8817 14815 8846 14818
rect 8817 14798 8823 14815
rect 8840 14814 8846 14815
rect 8931 14814 8934 14820
rect 8840 14800 8934 14814
rect 8840 14798 8846 14800
rect 8817 14795 8846 14798
rect 8931 14794 8934 14800
rect 8960 14794 8963 14820
rect 8977 14794 8980 14820
rect 9006 14814 9009 14820
rect 10173 14814 10176 14820
rect 9006 14800 10176 14814
rect 9006 14794 9009 14800
rect 10173 14794 10176 14800
rect 10202 14794 10205 14820
rect 10231 14815 10260 14818
rect 10231 14814 10237 14815
rect 10228 14798 10237 14814
rect 10254 14798 10260 14815
rect 10387 14815 10416 14818
rect 10228 14795 10260 14798
rect 10335 14805 10364 14808
rect 8701 14780 8704 14786
rect 8388 14766 8704 14780
rect 8701 14760 8704 14766
rect 8730 14780 8733 14786
rect 8885 14784 8888 14786
rect 8863 14781 8888 14784
rect 8863 14780 8869 14781
rect 8730 14766 8869 14780
rect 8730 14760 8733 14766
rect 8863 14764 8869 14766
rect 8886 14764 8888 14781
rect 8863 14761 8888 14764
rect 8885 14760 8888 14761
rect 8914 14760 8917 14786
rect 9691 14781 9720 14784
rect 9691 14764 9697 14781
rect 9714 14780 9720 14781
rect 10228 14780 10242 14795
rect 10335 14788 10341 14805
rect 10358 14788 10364 14805
rect 10387 14798 10393 14815
rect 10410 14798 10416 14815
rect 10435 14804 10441 14821
rect 10458 14804 10464 14821
rect 10435 14801 10464 14804
rect 10486 14815 10515 14818
rect 10387 14795 10416 14798
rect 10486 14798 10492 14815
rect 10509 14814 10515 14815
rect 10734 14814 10748 14902
rect 12059 14896 12062 14902
rect 12088 14896 12091 14922
rect 12565 14896 12568 14922
rect 12594 14916 12597 14922
rect 13025 14916 13028 14922
rect 12594 14902 13028 14916
rect 12594 14896 12597 14902
rect 13025 14896 13028 14902
rect 13054 14896 13057 14922
rect 15211 14917 15240 14920
rect 15211 14900 15217 14917
rect 15234 14916 15240 14917
rect 15785 14916 15788 14922
rect 15234 14902 15788 14916
rect 15234 14900 15240 14902
rect 15211 14897 15240 14900
rect 15785 14896 15788 14902
rect 15814 14896 15817 14922
rect 16108 14917 16137 14920
rect 16108 14900 16114 14917
rect 16131 14916 16137 14917
rect 16567 14916 16570 14922
rect 16131 14902 16570 14916
rect 16131 14900 16137 14902
rect 16108 14897 16137 14900
rect 16567 14896 16570 14902
rect 16596 14896 16599 14922
rect 12289 14862 12292 14888
rect 12318 14882 12321 14888
rect 12318 14868 13615 14882
rect 12318 14862 12321 14868
rect 10771 14828 10774 14854
rect 10800 14848 10803 14854
rect 11415 14848 11418 14854
rect 10800 14834 11418 14848
rect 10800 14828 10803 14834
rect 11415 14828 11418 14834
rect 11444 14828 11447 14854
rect 13601 14824 13615 14868
rect 13669 14862 13672 14888
rect 13698 14862 13701 14888
rect 13593 14821 13622 14824
rect 10509 14800 10748 14814
rect 11577 14815 11606 14818
rect 10509 14798 10515 14800
rect 10486 14795 10515 14798
rect 11577 14798 11583 14815
rect 11600 14814 11606 14815
rect 11691 14814 11694 14820
rect 11600 14800 11694 14814
rect 11600 14798 11606 14800
rect 11577 14795 11606 14798
rect 10335 14785 10364 14788
rect 9714 14766 10242 14780
rect 9714 14764 9720 14766
rect 9691 14761 9720 14764
rect 10343 14752 10357 14785
rect 10395 14780 10409 14795
rect 11691 14794 11694 14800
rect 11720 14794 11723 14820
rect 11737 14794 11740 14820
rect 11766 14814 11769 14820
rect 12289 14814 12292 14820
rect 11766 14800 12292 14814
rect 11766 14794 11769 14800
rect 12289 14794 12292 14800
rect 12318 14794 12321 14820
rect 13393 14794 13396 14820
rect 13422 14794 13425 14820
rect 13451 14815 13480 14818
rect 13451 14814 13457 14815
rect 13448 14798 13457 14814
rect 13474 14798 13480 14815
rect 13448 14795 13480 14798
rect 10541 14780 10544 14786
rect 10395 14766 10544 14780
rect 10541 14760 10544 14766
rect 10570 14760 10573 14786
rect 11627 14781 11656 14784
rect 11627 14764 11633 14781
rect 11650 14780 11656 14781
rect 11746 14780 11760 14794
rect 11650 14766 11760 14780
rect 12451 14781 12480 14784
rect 11650 14764 11656 14766
rect 11627 14761 11656 14764
rect 12451 14764 12457 14781
rect 12474 14780 12480 14781
rect 13448 14780 13462 14795
rect 13531 14794 13534 14820
rect 13560 14816 13563 14820
rect 13560 14813 13574 14816
rect 13568 14796 13574 14813
rect 13593 14804 13599 14821
rect 13616 14804 13622 14821
rect 13678 14818 13692 14862
rect 13807 14828 13810 14854
rect 13836 14848 13839 14854
rect 14175 14848 14178 14854
rect 13836 14834 14178 14848
rect 13836 14828 13839 14834
rect 14175 14828 14178 14834
rect 14204 14828 14207 14854
rect 16015 14828 16018 14854
rect 16044 14848 16047 14854
rect 16154 14849 16183 14852
rect 16154 14848 16160 14849
rect 16044 14834 16160 14848
rect 16044 14828 16047 14834
rect 16154 14832 16160 14834
rect 16177 14832 16183 14849
rect 16154 14829 16183 14832
rect 24157 14828 24160 14854
rect 24186 14848 24189 14854
rect 24341 14848 24344 14854
rect 24186 14834 24344 14848
rect 24186 14828 24189 14834
rect 24341 14828 24344 14834
rect 24370 14848 24373 14854
rect 24618 14849 24647 14852
rect 24618 14848 24624 14849
rect 24370 14834 24624 14848
rect 24370 14828 24373 14834
rect 24618 14832 24624 14834
rect 24641 14832 24647 14849
rect 24618 14829 24647 14832
rect 13715 14818 13718 14820
rect 13593 14801 13622 14804
rect 13655 14815 13692 14818
rect 13560 14794 13574 14796
rect 13655 14798 13661 14815
rect 13678 14800 13692 14815
rect 13706 14815 13718 14818
rect 13678 14798 13684 14800
rect 13655 14795 13684 14798
rect 13706 14798 13712 14815
rect 13706 14795 13718 14798
rect 13715 14794 13718 14795
rect 13744 14794 13747 14820
rect 15877 14794 15880 14820
rect 15906 14814 15909 14820
rect 15970 14815 15999 14818
rect 15970 14814 15976 14815
rect 15906 14800 15976 14814
rect 15906 14794 15909 14800
rect 15970 14798 15976 14800
rect 15993 14798 15999 14815
rect 15970 14795 15999 14798
rect 21535 14794 21538 14820
rect 21564 14814 21567 14820
rect 22041 14814 22044 14820
rect 21564 14800 22044 14814
rect 21564 14794 21567 14800
rect 22041 14794 22044 14800
rect 22070 14794 22073 14820
rect 24387 14794 24390 14820
rect 24416 14814 24419 14820
rect 24755 14814 24758 14820
rect 24784 14818 24787 14820
rect 24784 14815 24802 14818
rect 24416 14800 24758 14814
rect 24416 14794 24419 14800
rect 24755 14794 24758 14800
rect 24796 14798 24802 14815
rect 24784 14795 24802 14798
rect 24784 14794 24787 14795
rect 13545 14793 13574 14794
rect 12474 14766 13462 14780
rect 12474 14764 12480 14766
rect 12451 14761 12480 14764
rect 13807 14760 13810 14786
rect 13836 14780 13839 14786
rect 13945 14780 13948 14786
rect 13836 14766 13948 14780
rect 13836 14760 13839 14766
rect 13945 14760 13948 14766
rect 13974 14780 13977 14786
rect 14221 14780 14224 14786
rect 13974 14766 14224 14780
rect 13974 14760 13977 14766
rect 14221 14760 14224 14766
rect 14250 14780 14253 14786
rect 14405 14784 14408 14786
rect 14336 14781 14365 14784
rect 14336 14780 14342 14781
rect 14250 14766 14342 14780
rect 14250 14760 14253 14766
rect 14336 14764 14342 14766
rect 14359 14764 14365 14781
rect 14336 14761 14365 14764
rect 14387 14781 14408 14784
rect 14387 14764 14393 14781
rect 14387 14761 14408 14764
rect 14405 14760 14408 14761
rect 14434 14760 14437 14786
rect 16016 14781 16045 14784
rect 16016 14764 16022 14781
rect 16039 14780 16045 14781
rect 16153 14780 16156 14786
rect 16039 14766 16156 14780
rect 16039 14764 16045 14766
rect 16016 14761 16045 14764
rect 16153 14760 16156 14766
rect 16182 14760 16185 14786
rect 22050 14780 22064 14794
rect 24825 14781 24854 14784
rect 24825 14780 24831 14781
rect 22050 14766 24831 14780
rect 24825 14764 24831 14766
rect 24848 14764 24854 14781
rect 24825 14761 24854 14764
rect 3181 14726 3184 14752
rect 3210 14726 3213 14752
rect 4838 14747 4867 14750
rect 4838 14730 4844 14747
rect 4861 14746 4867 14747
rect 5941 14746 5944 14752
rect 4861 14732 5944 14746
rect 4861 14730 4867 14732
rect 4838 14727 4867 14730
rect 5941 14726 5944 14732
rect 5970 14726 5973 14752
rect 10173 14726 10176 14752
rect 10202 14726 10205 14752
rect 10343 14732 10360 14752
rect 10357 14726 10360 14732
rect 10386 14726 10389 14752
rect 13624 14747 13653 14750
rect 13624 14730 13630 14747
rect 13647 14746 13653 14747
rect 13899 14746 13902 14752
rect 13647 14732 13902 14746
rect 13647 14730 13653 14732
rect 13624 14727 13653 14730
rect 13899 14726 13902 14732
rect 13928 14726 13931 14752
rect 16061 14726 16064 14752
rect 16090 14726 16093 14752
rect 25653 14747 25682 14750
rect 25653 14730 25659 14747
rect 25676 14746 25682 14747
rect 25905 14746 25908 14752
rect 25676 14732 25908 14746
rect 25676 14730 25682 14732
rect 25653 14727 25682 14730
rect 25905 14726 25908 14732
rect 25934 14726 25937 14752
rect 3036 14664 29992 14712
rect 4815 14645 4844 14648
rect 4815 14628 4821 14645
rect 4838 14644 4844 14645
rect 4929 14644 4932 14650
rect 4838 14630 4932 14644
rect 4838 14628 4844 14630
rect 4815 14625 4844 14628
rect 4929 14624 4932 14630
rect 4958 14624 4961 14650
rect 7459 14624 7462 14650
rect 7488 14644 7491 14650
rect 7713 14645 7742 14648
rect 7713 14644 7719 14645
rect 7488 14630 7719 14644
rect 7488 14624 7491 14630
rect 7713 14628 7719 14630
rect 7736 14628 7742 14645
rect 7713 14625 7742 14628
rect 11691 14624 11694 14650
rect 11720 14644 11723 14650
rect 13417 14645 13446 14648
rect 11720 14630 11806 14644
rect 11720 14624 11723 14630
rect 3825 14590 3828 14616
rect 3854 14610 3857 14616
rect 9345 14614 9348 14616
rect 3979 14611 4008 14614
rect 3979 14610 3985 14611
rect 3854 14596 3985 14610
rect 3854 14590 3857 14596
rect 3979 14594 3985 14596
rect 4002 14594 4008 14611
rect 3979 14591 4008 14594
rect 6889 14611 6918 14614
rect 6889 14594 6895 14611
rect 6912 14610 6918 14611
rect 9327 14611 9348 14614
rect 6912 14596 7022 14610
rect 6912 14594 6918 14596
rect 6889 14591 6918 14594
rect 3181 14556 3184 14582
rect 3210 14576 3213 14582
rect 3411 14576 3414 14582
rect 3210 14562 3414 14576
rect 3210 14556 3213 14562
rect 3411 14556 3414 14562
rect 3440 14576 3443 14582
rect 3935 14577 3964 14580
rect 3935 14576 3941 14577
rect 3440 14562 3941 14576
rect 3440 14556 3443 14562
rect 3935 14560 3941 14562
rect 3958 14560 3964 14577
rect 3935 14557 3964 14560
rect 5895 14556 5898 14582
rect 5924 14576 5927 14582
rect 5924 14562 6217 14576
rect 5924 14556 5927 14562
rect 3319 14522 3322 14548
rect 3348 14542 3351 14548
rect 3780 14543 3809 14546
rect 3780 14542 3786 14543
rect 3348 14528 3786 14542
rect 3348 14522 3351 14528
rect 3780 14526 3786 14528
rect 3803 14526 3809 14543
rect 6203 14542 6217 14562
rect 6815 14556 6818 14582
rect 6844 14580 6847 14582
rect 6844 14577 6862 14580
rect 6856 14560 6862 14577
rect 7008 14576 7022 14596
rect 9327 14594 9333 14611
rect 9327 14591 9348 14594
rect 9345 14590 9348 14591
rect 9374 14590 9377 14616
rect 10265 14590 10268 14616
rect 10294 14610 10297 14616
rect 11737 14610 11740 14616
rect 10294 14596 11740 14610
rect 10294 14590 10297 14596
rect 11737 14590 11740 14596
rect 11766 14590 11769 14616
rect 11792 14610 11806 14630
rect 13417 14628 13423 14645
rect 13440 14644 13446 14645
rect 13531 14644 13534 14650
rect 13440 14630 13534 14644
rect 13440 14628 13446 14630
rect 13417 14625 13446 14628
rect 13531 14624 13534 14630
rect 13560 14624 13563 14650
rect 12593 14611 12622 14614
rect 11792 14596 12542 14610
rect 12528 14582 12542 14596
rect 12593 14594 12599 14611
rect 12616 14610 12622 14611
rect 12657 14610 12660 14616
rect 12616 14596 12660 14610
rect 12616 14594 12622 14596
rect 12593 14591 12622 14594
rect 12657 14590 12660 14596
rect 12686 14590 12689 14616
rect 15417 14614 15420 14616
rect 15399 14611 15420 14614
rect 15399 14594 15405 14611
rect 15399 14591 15420 14594
rect 15417 14590 15420 14591
rect 15446 14590 15449 14616
rect 26393 14611 26422 14614
rect 26393 14594 26399 14611
rect 26416 14610 26422 14611
rect 26457 14610 26460 14616
rect 26416 14596 26460 14610
rect 26416 14594 26422 14596
rect 26393 14591 26422 14594
rect 26457 14590 26460 14596
rect 26486 14590 26489 14616
rect 7091 14576 7094 14582
rect 7008 14562 7094 14576
rect 6844 14557 6862 14560
rect 6844 14556 6847 14557
rect 7091 14556 7094 14562
rect 7120 14556 7123 14582
rect 8931 14556 8934 14582
rect 8960 14576 8963 14582
rect 9253 14576 9256 14582
rect 9282 14580 9285 14582
rect 9282 14577 9300 14580
rect 8960 14562 9256 14576
rect 8960 14556 8963 14562
rect 9253 14556 9256 14562
rect 9294 14560 9300 14577
rect 9282 14557 9300 14560
rect 9282 14556 9285 14557
rect 11415 14556 11418 14582
rect 11444 14576 11447 14582
rect 12381 14576 12384 14582
rect 11444 14562 12384 14576
rect 11444 14556 11447 14562
rect 12381 14556 12384 14562
rect 12410 14556 12413 14582
rect 12519 14556 12522 14582
rect 12548 14580 12551 14582
rect 12548 14577 12566 14580
rect 12560 14560 12566 14577
rect 12548 14557 12566 14560
rect 12548 14556 12551 14557
rect 14221 14556 14224 14582
rect 14250 14576 14253 14582
rect 15343 14577 15372 14580
rect 15343 14576 15349 14577
rect 14250 14562 15349 14576
rect 14250 14556 14253 14562
rect 15343 14560 15349 14562
rect 15366 14576 15372 14577
rect 15463 14576 15466 14582
rect 15366 14562 15466 14576
rect 15366 14560 15372 14562
rect 15343 14557 15372 14560
rect 15463 14556 15466 14562
rect 15492 14556 15495 14582
rect 26135 14556 26138 14582
rect 26164 14576 26167 14582
rect 26343 14577 26372 14580
rect 26343 14576 26349 14577
rect 26164 14562 26349 14576
rect 26164 14556 26167 14562
rect 26343 14560 26349 14562
rect 26366 14576 26372 14577
rect 28297 14576 28300 14582
rect 26366 14562 28300 14576
rect 26366 14560 26372 14562
rect 26343 14557 26372 14560
rect 28297 14556 28300 14562
rect 28326 14556 28329 14582
rect 29355 14556 29358 14582
rect 29384 14556 29387 14582
rect 29447 14556 29450 14582
rect 29476 14556 29479 14582
rect 6678 14543 6707 14546
rect 6678 14542 6684 14543
rect 6203 14528 6684 14542
rect 3780 14523 3809 14526
rect 6678 14526 6684 14528
rect 6701 14526 6707 14543
rect 6678 14523 6707 14526
rect 6686 14474 6700 14523
rect 8517 14522 8520 14548
rect 8546 14542 8549 14548
rect 9115 14542 9118 14548
rect 8546 14528 9118 14542
rect 8546 14522 8549 14528
rect 9115 14522 9118 14528
rect 9144 14522 9147 14548
rect 14175 14522 14178 14548
rect 14204 14542 14207 14548
rect 15187 14542 15190 14548
rect 14204 14528 15190 14542
rect 14204 14522 14207 14528
rect 15187 14522 15190 14528
rect 15216 14522 15219 14548
rect 25997 14522 26000 14548
rect 26026 14542 26029 14548
rect 26182 14543 26211 14546
rect 26182 14542 26188 14543
rect 26026 14528 26188 14542
rect 26026 14522 26029 14528
rect 26182 14526 26188 14528
rect 26205 14526 26211 14543
rect 26182 14523 26211 14526
rect 6861 14474 6864 14480
rect 6686 14460 6864 14474
rect 6861 14454 6864 14460
rect 6890 14474 6893 14480
rect 7275 14474 7278 14480
rect 6890 14460 7278 14474
rect 6890 14454 6893 14460
rect 7275 14454 7278 14460
rect 7304 14454 7307 14480
rect 10151 14475 10180 14478
rect 10151 14458 10157 14475
rect 10174 14474 10180 14475
rect 10357 14474 10360 14480
rect 10174 14460 10360 14474
rect 10174 14458 10180 14460
rect 10151 14455 10180 14458
rect 10357 14454 10360 14460
rect 10386 14454 10389 14480
rect 16199 14454 16202 14480
rect 16228 14478 16231 14480
rect 16228 14475 16252 14478
rect 16228 14458 16229 14475
rect 16246 14458 16252 14475
rect 16228 14455 16252 14458
rect 16228 14454 16231 14455
rect 22915 14454 22918 14480
rect 22944 14474 22947 14480
rect 24295 14474 24298 14480
rect 22944 14460 24298 14474
rect 22944 14454 22947 14460
rect 24295 14454 24298 14460
rect 24324 14454 24327 14480
rect 27217 14475 27246 14478
rect 27217 14458 27223 14475
rect 27240 14474 27246 14475
rect 27515 14474 27518 14480
rect 27240 14460 27518 14474
rect 27240 14458 27246 14460
rect 27217 14455 27246 14458
rect 27515 14454 27518 14460
rect 27544 14454 27547 14480
rect 29402 14475 29431 14478
rect 29402 14458 29408 14475
rect 29425 14474 29431 14475
rect 29585 14474 29588 14480
rect 29425 14460 29588 14474
rect 29425 14458 29431 14460
rect 29402 14455 29431 14458
rect 29585 14454 29588 14460
rect 29614 14454 29617 14480
rect 3036 14392 29992 14440
rect 3319 14372 3322 14378
rect 3144 14358 3322 14372
rect 3144 14308 3158 14358
rect 3319 14352 3322 14358
rect 3348 14352 3351 14378
rect 4171 14373 4200 14376
rect 4171 14356 4177 14373
rect 4194 14372 4200 14373
rect 4975 14372 4978 14378
rect 4194 14358 4978 14372
rect 4194 14356 4200 14358
rect 4171 14353 4200 14356
rect 4975 14352 4978 14358
rect 5004 14352 5007 14378
rect 6793 14373 6822 14376
rect 6793 14356 6799 14373
rect 6816 14372 6822 14373
rect 6907 14372 6910 14378
rect 6816 14358 6910 14372
rect 6816 14356 6822 14358
rect 6793 14353 6822 14356
rect 6907 14352 6910 14358
rect 6936 14352 6939 14378
rect 8679 14373 8708 14376
rect 8679 14356 8685 14373
rect 8702 14372 8708 14373
rect 8839 14372 8842 14378
rect 8702 14358 8842 14372
rect 8702 14356 8708 14358
rect 8679 14353 8708 14356
rect 8839 14352 8842 14358
rect 8868 14352 8871 14378
rect 14291 14373 14320 14376
rect 13218 14358 14106 14372
rect 3136 14305 3165 14308
rect 3136 14288 3142 14305
rect 3159 14288 3165 14305
rect 3136 14285 3165 14288
rect 4975 14284 4978 14310
rect 5004 14304 5007 14310
rect 5251 14304 5254 14310
rect 5004 14290 5254 14304
rect 5004 14284 5007 14290
rect 5251 14284 5254 14290
rect 5280 14284 5283 14310
rect 5711 14284 5714 14310
rect 5740 14304 5743 14310
rect 5758 14305 5787 14308
rect 5758 14304 5764 14305
rect 5740 14290 5764 14304
rect 5740 14284 5743 14290
rect 5758 14288 5764 14290
rect 5781 14288 5787 14305
rect 5758 14285 5787 14288
rect 7275 14284 7278 14310
rect 7304 14304 7307 14310
rect 7643 14304 7646 14310
rect 7304 14290 7646 14304
rect 7304 14284 7307 14290
rect 7643 14284 7646 14290
rect 7672 14284 7675 14310
rect 11899 14305 11928 14308
rect 11899 14288 11905 14305
rect 11922 14304 11928 14305
rect 11922 14290 12358 14304
rect 11922 14288 11928 14290
rect 11899 14285 11928 14288
rect 3181 14250 3184 14276
rect 3210 14270 3213 14276
rect 3291 14271 3320 14274
rect 3291 14270 3297 14271
rect 3210 14256 3297 14270
rect 3210 14250 3213 14256
rect 3291 14254 3297 14256
rect 3314 14254 3320 14271
rect 3457 14270 3460 14276
rect 3291 14251 3320 14254
rect 3443 14250 3460 14270
rect 3486 14250 3489 14276
rect 4791 14250 4794 14276
rect 4820 14270 4823 14276
rect 5113 14270 5116 14276
rect 4820 14256 5116 14270
rect 4820 14250 4823 14256
rect 5113 14250 5116 14256
rect 5142 14270 5145 14276
rect 5919 14271 5948 14274
rect 5919 14270 5925 14271
rect 5142 14256 5925 14270
rect 5142 14250 5145 14256
rect 5919 14254 5925 14256
rect 5942 14270 5948 14271
rect 6033 14270 6036 14276
rect 5942 14256 6036 14270
rect 5942 14254 5948 14256
rect 5919 14251 5948 14254
rect 6033 14250 6036 14256
rect 6062 14250 6065 14276
rect 6953 14270 6956 14276
rect 6088 14256 6956 14270
rect 3347 14237 3376 14240
rect 3347 14220 3353 14237
rect 3370 14236 3376 14237
rect 3443 14236 3457 14250
rect 3370 14222 3457 14236
rect 5969 14237 5998 14240
rect 3370 14220 3376 14222
rect 3347 14217 3376 14220
rect 5969 14220 5975 14237
rect 5992 14236 5998 14237
rect 6088 14236 6102 14256
rect 6953 14250 6956 14256
rect 6982 14250 6985 14276
rect 7781 14250 7784 14276
rect 7810 14274 7813 14276
rect 7810 14271 7828 14274
rect 7822 14254 7828 14271
rect 7810 14251 7828 14254
rect 7843 14271 7872 14274
rect 7843 14254 7849 14271
rect 7866 14270 7872 14271
rect 8701 14270 8704 14276
rect 7866 14256 8704 14270
rect 7866 14254 7872 14256
rect 7843 14251 7872 14254
rect 7810 14250 7813 14251
rect 8701 14250 8704 14256
rect 8730 14250 8733 14276
rect 10771 14250 10774 14276
rect 10800 14270 10803 14276
rect 10864 14271 10893 14274
rect 10864 14270 10870 14271
rect 10800 14256 10870 14270
rect 10800 14250 10803 14256
rect 10864 14254 10870 14256
rect 10887 14254 10893 14271
rect 10864 14251 10893 14254
rect 11001 14250 11004 14276
rect 11030 14274 11033 14276
rect 11030 14271 11054 14274
rect 11030 14254 11031 14271
rect 11048 14270 11054 14271
rect 11139 14270 11142 14276
rect 11048 14256 11142 14270
rect 11048 14254 11054 14256
rect 11030 14251 11054 14254
rect 11030 14250 11033 14251
rect 11139 14250 11142 14256
rect 11168 14250 11171 14276
rect 12151 14250 12154 14276
rect 12180 14250 12183 14276
rect 12197 14250 12200 14276
rect 12226 14250 12229 14276
rect 12344 14274 12358 14290
rect 12336 14271 12365 14274
rect 12336 14254 12342 14271
rect 12359 14254 12365 14271
rect 12336 14251 12365 14254
rect 12381 14250 12384 14276
rect 12410 14270 12413 14276
rect 13218 14270 13232 14358
rect 14092 14338 14106 14358
rect 14291 14356 14297 14373
rect 14314 14372 14320 14373
rect 14497 14372 14500 14378
rect 14314 14358 14500 14372
rect 14314 14356 14320 14358
rect 14291 14353 14320 14356
rect 14497 14352 14500 14358
rect 14526 14352 14529 14378
rect 15141 14352 15144 14378
rect 15170 14372 15173 14378
rect 17165 14372 17168 14378
rect 15170 14358 17168 14372
rect 15170 14352 15173 14358
rect 17165 14352 17168 14358
rect 17194 14352 17197 14378
rect 22685 14352 22688 14378
rect 22714 14372 22717 14378
rect 28251 14372 28254 14378
rect 22714 14358 25974 14372
rect 22714 14352 22717 14358
rect 15647 14338 15650 14344
rect 14092 14324 15650 14338
rect 15647 14318 15650 14324
rect 15676 14318 15679 14344
rect 21489 14318 21492 14344
rect 21518 14338 21521 14344
rect 22870 14339 22899 14342
rect 22870 14338 22876 14339
rect 21518 14324 22876 14338
rect 21518 14318 21521 14324
rect 22870 14322 22876 14324
rect 22893 14322 22899 14339
rect 22870 14319 22899 14322
rect 25813 14318 25816 14344
rect 25842 14318 25845 14344
rect 25905 14318 25908 14344
rect 25934 14318 25937 14344
rect 17304 14305 17333 14308
rect 17304 14288 17310 14305
rect 17327 14304 17333 14305
rect 17764 14305 17793 14308
rect 17327 14290 17740 14304
rect 17327 14288 17333 14290
rect 17304 14285 17333 14288
rect 12410 14256 13232 14270
rect 12410 14250 12413 14256
rect 13255 14250 13258 14276
rect 13284 14250 13287 14276
rect 13455 14271 13484 14274
rect 13455 14270 13461 14271
rect 13310 14256 13461 14270
rect 11093 14240 11096 14242
rect 5992 14222 6102 14236
rect 11075 14237 11096 14240
rect 5992 14220 5998 14222
rect 5969 14217 5998 14220
rect 11075 14220 11081 14237
rect 11075 14217 11096 14220
rect 11093 14216 11096 14217
rect 11122 14216 11125 14242
rect 12289 14216 12292 14242
rect 12318 14216 12321 14242
rect 12243 14182 12246 14208
rect 12272 14182 12275 14208
rect 12335 14182 12338 14208
rect 12364 14202 12367 14208
rect 13310 14202 13324 14256
rect 13455 14254 13461 14256
rect 13478 14254 13484 14271
rect 13807 14270 13810 14276
rect 13455 14251 13484 14254
rect 13586 14256 13810 14270
rect 13416 14237 13445 14240
rect 13416 14220 13422 14237
rect 13439 14236 13445 14237
rect 13586 14236 13600 14256
rect 13807 14250 13810 14256
rect 13836 14250 13839 14276
rect 17671 14250 17674 14276
rect 17700 14250 17703 14276
rect 17726 14270 17740 14290
rect 17764 14288 17770 14305
rect 17787 14304 17793 14305
rect 17901 14304 17904 14310
rect 17787 14290 17904 14304
rect 17787 14288 17793 14290
rect 17764 14285 17793 14288
rect 17901 14284 17904 14290
rect 17930 14284 17933 14310
rect 19281 14284 19284 14310
rect 19310 14304 19313 14310
rect 21214 14305 21243 14308
rect 21214 14304 21220 14305
rect 19310 14290 21220 14304
rect 19310 14284 19313 14290
rect 21214 14288 21220 14290
rect 21237 14288 21243 14305
rect 21214 14285 21243 14288
rect 21351 14284 21354 14310
rect 21380 14284 21383 14310
rect 24341 14284 24344 14310
rect 24370 14284 24373 14310
rect 25377 14305 25406 14308
rect 25377 14288 25383 14305
rect 25400 14304 25406 14305
rect 25822 14304 25836 14318
rect 25400 14290 25709 14304
rect 25822 14290 25851 14304
rect 25400 14288 25406 14290
rect 25377 14285 25406 14288
rect 17856 14271 17885 14274
rect 17856 14270 17862 14271
rect 17726 14256 17862 14270
rect 17772 14242 17786 14256
rect 17856 14254 17862 14256
rect 17879 14254 17885 14271
rect 17856 14251 17885 14254
rect 19373 14250 19376 14276
rect 19402 14270 19405 14276
rect 19512 14271 19541 14274
rect 19512 14270 19518 14271
rect 19402 14256 19518 14270
rect 19402 14250 19405 14256
rect 19512 14254 19518 14256
rect 19535 14254 19541 14271
rect 19512 14251 19541 14254
rect 19879 14250 19882 14276
rect 19908 14270 19911 14276
rect 19926 14271 19955 14274
rect 19926 14270 19932 14271
rect 19908 14256 19932 14270
rect 19908 14250 19911 14256
rect 19926 14254 19932 14256
rect 19949 14254 19955 14271
rect 19926 14251 19955 14254
rect 21121 14250 21124 14276
rect 21150 14270 21153 14276
rect 21260 14271 21289 14274
rect 21260 14270 21266 14271
rect 21150 14256 21266 14270
rect 21150 14250 21153 14256
rect 21260 14254 21266 14256
rect 21283 14254 21289 14271
rect 21260 14251 21289 14254
rect 22869 14250 22872 14276
rect 22898 14250 22901 14276
rect 23008 14271 23037 14274
rect 23008 14254 23014 14271
rect 23031 14270 23037 14271
rect 24663 14270 24666 14276
rect 23031 14256 24666 14270
rect 23031 14254 23037 14256
rect 23008 14251 23037 14254
rect 24663 14250 24666 14256
rect 24692 14250 24695 14276
rect 25629 14250 25632 14276
rect 25658 14250 25661 14276
rect 25695 14274 25709 14290
rect 25687 14271 25716 14274
rect 25687 14254 25693 14271
rect 25710 14254 25716 14271
rect 25687 14251 25716 14254
rect 25767 14250 25770 14276
rect 25796 14274 25799 14276
rect 25837 14274 25851 14290
rect 25914 14275 25928 14318
rect 25960 14304 25974 14358
rect 25796 14271 25810 14274
rect 25804 14254 25810 14271
rect 25796 14251 25810 14254
rect 25829 14271 25858 14274
rect 25899 14272 25928 14275
rect 25950 14290 25974 14304
rect 27708 14358 28254 14372
rect 27708 14304 27722 14358
rect 28251 14352 28254 14358
rect 28280 14352 28283 14378
rect 27708 14290 27768 14304
rect 25950 14274 25964 14290
rect 25829 14254 25835 14271
rect 25852 14254 25858 14271
rect 25829 14251 25858 14254
rect 25884 14269 25928 14272
rect 25884 14252 25890 14269
rect 25907 14261 25928 14269
rect 25942 14271 25971 14274
rect 25907 14252 25913 14261
rect 25796 14250 25799 14251
rect 25884 14249 25913 14252
rect 25942 14254 25948 14271
rect 25965 14254 25971 14271
rect 25942 14251 25971 14254
rect 25997 14250 26000 14276
rect 26026 14270 26029 14276
rect 27699 14270 27702 14276
rect 26026 14256 27702 14270
rect 26026 14250 26029 14256
rect 27699 14250 27702 14256
rect 27728 14250 27731 14276
rect 27754 14270 27768 14290
rect 27855 14271 27884 14274
rect 27855 14270 27861 14271
rect 27754 14256 27861 14270
rect 27855 14254 27861 14256
rect 27878 14254 27884 14271
rect 28343 14270 28346 14276
rect 27855 14251 27884 14254
rect 28030 14256 28346 14270
rect 13439 14222 13600 14236
rect 13439 14220 13445 14222
rect 13416 14217 13445 14220
rect 17763 14216 17766 14242
rect 17792 14216 17795 14242
rect 19696 14237 19725 14240
rect 19696 14220 19702 14237
rect 19719 14236 19725 14237
rect 22962 14237 22991 14240
rect 22962 14236 22968 14237
rect 19719 14222 22968 14236
rect 19719 14220 19725 14222
rect 19696 14217 19725 14220
rect 22962 14220 22968 14222
rect 22985 14236 22991 14237
rect 23099 14236 23102 14242
rect 22985 14222 23102 14236
rect 22985 14220 22991 14222
rect 22962 14217 22991 14220
rect 23099 14216 23102 14222
rect 23128 14216 23131 14242
rect 24387 14216 24390 14242
rect 24416 14236 24419 14242
rect 24571 14240 24574 14242
rect 24502 14237 24531 14240
rect 24502 14236 24508 14237
rect 24416 14222 24508 14236
rect 24416 14216 24419 14222
rect 24502 14220 24508 14222
rect 24525 14220 24531 14237
rect 24502 14217 24531 14220
rect 24553 14237 24574 14240
rect 24553 14220 24559 14237
rect 24553 14217 24574 14220
rect 24571 14216 24574 14217
rect 24600 14216 24603 14242
rect 27911 14237 27940 14240
rect 27911 14220 27917 14237
rect 27934 14236 27940 14237
rect 28030 14236 28044 14256
rect 28343 14250 28346 14256
rect 28372 14270 28375 14276
rect 28435 14270 28438 14276
rect 28372 14256 28438 14270
rect 28372 14250 28375 14256
rect 28435 14250 28438 14256
rect 28464 14250 28467 14276
rect 27934 14222 28044 14236
rect 27934 14220 27940 14222
rect 27911 14217 27940 14220
rect 12364 14188 13324 14202
rect 12364 14182 12367 14188
rect 17211 14182 17214 14208
rect 17240 14202 17243 14208
rect 17396 14203 17425 14206
rect 17396 14202 17402 14203
rect 17240 14188 17402 14202
rect 17240 14182 17243 14188
rect 17396 14186 17402 14188
rect 17419 14186 17425 14203
rect 17396 14183 17425 14186
rect 17717 14182 17720 14208
rect 17746 14182 17749 14208
rect 17809 14182 17812 14208
rect 17838 14182 17841 14208
rect 19511 14182 19514 14208
rect 19540 14182 19543 14208
rect 21352 14203 21381 14206
rect 21352 14186 21358 14203
rect 21375 14202 21381 14203
rect 21443 14202 21446 14208
rect 21375 14188 21446 14202
rect 21375 14186 21381 14188
rect 21352 14183 21381 14186
rect 21443 14182 21446 14188
rect 21472 14182 21475 14208
rect 25860 14203 25889 14206
rect 25860 14186 25866 14203
rect 25883 14202 25889 14203
rect 26825 14202 26828 14208
rect 25883 14188 26828 14202
rect 25883 14186 25889 14188
rect 25860 14183 25889 14186
rect 26825 14182 26828 14188
rect 26854 14182 26857 14208
rect 28573 14182 28576 14208
rect 28602 14202 28605 14208
rect 28735 14203 28764 14206
rect 28735 14202 28741 14203
rect 28602 14188 28741 14202
rect 28602 14182 28605 14188
rect 28735 14186 28741 14188
rect 28758 14186 28764 14203
rect 28735 14183 28764 14186
rect 3036 14120 29992 14168
rect 11093 14080 11096 14106
rect 11122 14100 11125 14106
rect 14451 14100 14454 14106
rect 11122 14086 14454 14100
rect 11122 14080 11125 14086
rect 14451 14080 14454 14086
rect 14480 14080 14483 14106
rect 17763 14080 17766 14106
rect 17792 14080 17795 14106
rect 19879 14080 19882 14106
rect 19908 14100 19911 14106
rect 19908 14086 20500 14100
rect 19908 14080 19911 14086
rect 3181 14046 3184 14072
rect 3210 14066 3213 14072
rect 4727 14067 4756 14070
rect 3210 14052 4699 14066
rect 3210 14046 3213 14052
rect 4685 14036 4699 14052
rect 4727 14050 4733 14067
rect 4750 14066 4756 14067
rect 6401 14066 6404 14072
rect 4750 14052 4862 14066
rect 4750 14050 4756 14052
rect 4727 14047 4756 14050
rect 4677 14033 4706 14036
rect 4677 14016 4683 14033
rect 4700 14032 4706 14033
rect 4791 14032 4794 14038
rect 4700 14018 4794 14032
rect 4700 14016 4706 14018
rect 4677 14013 4706 14016
rect 4791 14012 4794 14018
rect 4820 14012 4823 14038
rect 4848 14032 4862 14052
rect 6088 14052 6404 14066
rect 5251 14032 5254 14038
rect 4848 14018 5254 14032
rect 5251 14012 5254 14018
rect 5280 14012 5283 14038
rect 6088 14036 6102 14052
rect 6401 14046 6404 14052
rect 6430 14046 6433 14072
rect 9714 14067 9743 14070
rect 9714 14050 9720 14067
rect 9737 14066 9743 14067
rect 12289 14066 12292 14072
rect 9737 14052 12292 14066
rect 9737 14050 9743 14052
rect 9714 14047 9743 14050
rect 12289 14046 12292 14052
rect 12318 14046 12321 14072
rect 17257 14066 17260 14072
rect 15242 14052 17260 14066
rect 6080 14033 6109 14036
rect 6080 14016 6086 14033
rect 6103 14016 6109 14033
rect 6080 14013 6109 14016
rect 6127 14033 6156 14036
rect 6127 14016 6133 14033
rect 6150 14016 6156 14033
rect 6127 14013 6156 14016
rect 6218 14033 6247 14036
rect 6218 14016 6224 14033
rect 6241 14016 6247 14033
rect 6218 14013 6247 14016
rect 3319 13978 3322 14004
rect 3348 13998 3351 14004
rect 4516 13999 4545 14002
rect 4516 13998 4522 13999
rect 3348 13984 4522 13998
rect 3348 13978 3351 13984
rect 4516 13982 4522 13984
rect 4539 13982 4545 13999
rect 4516 13979 4545 13982
rect 5551 13999 5580 14002
rect 5551 13982 5557 13999
rect 5574 13998 5580 13999
rect 6134 13998 6148 14013
rect 5574 13984 6148 13998
rect 6226 13998 6240 14013
rect 6263 14012 6266 14038
rect 6292 14012 6295 14038
rect 6333 14033 6362 14036
rect 6333 14016 6339 14033
rect 6356 14032 6362 14033
rect 6447 14032 6450 14038
rect 6356 14018 6450 14032
rect 6356 14016 6362 14018
rect 6333 14013 6362 14016
rect 6447 14012 6450 14018
rect 6476 14032 6479 14038
rect 6476 14018 8402 14032
rect 6476 14012 6479 14018
rect 8388 13998 8402 14018
rect 9621 14012 9624 14038
rect 9650 14012 9653 14038
rect 9759 14012 9762 14038
rect 9788 14012 9791 14038
rect 9824 14033 9853 14036
rect 9824 14032 9830 14033
rect 9814 14016 9830 14032
rect 9847 14032 9853 14033
rect 9847 14018 11047 14032
rect 9847 14016 9853 14018
rect 9814 14013 9853 14016
rect 9814 13998 9828 14013
rect 6226 13984 6332 13998
rect 8388 13984 9828 13998
rect 5574 13982 5580 13984
rect 5551 13979 5580 13982
rect 4524 13930 4538 13979
rect 6318 13970 6332 13984
rect 6309 13944 6312 13970
rect 6338 13944 6341 13970
rect 11033 13964 11047 14018
rect 12298 13998 12312 14046
rect 15242 14036 15256 14052
rect 17257 14046 17260 14052
rect 17286 14046 17289 14072
rect 19373 14046 19376 14072
rect 19402 14066 19405 14072
rect 20486 14066 20500 14086
rect 20615 14080 20618 14106
rect 20644 14100 20647 14106
rect 21351 14100 21354 14106
rect 20644 14086 21354 14100
rect 20644 14080 20647 14086
rect 21351 14080 21354 14086
rect 21380 14080 21383 14106
rect 21443 14080 21446 14106
rect 21472 14080 21475 14106
rect 22823 14080 22826 14106
rect 22852 14100 22855 14106
rect 24111 14100 24114 14106
rect 22852 14086 24114 14100
rect 22852 14080 22855 14086
rect 24111 14080 24114 14086
rect 24140 14100 24143 14106
rect 25813 14100 25816 14106
rect 24140 14086 25816 14100
rect 24140 14080 24143 14086
rect 25813 14080 25816 14086
rect 25842 14080 25845 14106
rect 27423 14100 27426 14106
rect 27294 14086 27426 14100
rect 21489 14066 21492 14072
rect 19402 14052 19948 14066
rect 20486 14052 20546 14066
rect 19402 14046 19405 14052
rect 15234 14033 15263 14036
rect 15234 14016 15240 14033
rect 15257 14016 15263 14033
rect 15234 14013 15263 14016
rect 15280 14033 15309 14036
rect 15280 14016 15286 14033
rect 15303 14032 15309 14033
rect 15325 14032 15328 14038
rect 15303 14018 15328 14032
rect 15303 14016 15309 14018
rect 15280 14013 15309 14016
rect 15325 14012 15328 14018
rect 15354 14012 15357 14038
rect 15372 14033 15401 14036
rect 15372 14016 15378 14033
rect 15395 14016 15401 14033
rect 15372 14013 15401 14016
rect 15187 13998 15190 14004
rect 12298 13984 15190 13998
rect 15187 13978 15190 13984
rect 15216 13998 15219 14004
rect 15380 13998 15394 14013
rect 15417 14012 15420 14038
rect 15446 14012 15449 14038
rect 15464 14033 15493 14036
rect 15464 14016 15470 14033
rect 15487 14032 15493 14033
rect 15647 14032 15650 14038
rect 15487 14018 15650 14032
rect 15487 14016 15493 14018
rect 15464 14013 15493 14016
rect 15647 14012 15650 14018
rect 15676 14012 15679 14038
rect 16751 14012 16754 14038
rect 16780 14032 16783 14038
rect 17202 14033 17231 14036
rect 17202 14032 17208 14033
rect 16780 14018 17208 14032
rect 16780 14012 16783 14018
rect 17202 14016 17208 14018
rect 17225 14016 17231 14033
rect 17202 14013 17231 14016
rect 17671 14012 17674 14038
rect 17700 14032 17703 14038
rect 19879 14032 19882 14038
rect 17700 14018 19882 14032
rect 17700 14012 17703 14018
rect 19879 14012 19882 14018
rect 19908 14012 19911 14038
rect 19934 14032 19948 14052
rect 19971 14032 19974 14038
rect 19934 14018 19974 14032
rect 19971 14012 19974 14018
rect 20000 14032 20003 14038
rect 20532 14036 20546 14052
rect 21360 14052 21492 14066
rect 21360 14036 21374 14052
rect 21489 14046 21492 14052
rect 21518 14046 21521 14072
rect 26181 14070 26184 14072
rect 26163 14067 26184 14070
rect 26163 14050 26169 14067
rect 26163 14047 26184 14050
rect 26181 14046 26184 14047
rect 26210 14046 26213 14072
rect 20294 14033 20323 14036
rect 20294 14032 20300 14033
rect 20000 14018 20300 14032
rect 20000 14012 20003 14018
rect 20294 14016 20300 14018
rect 20317 14016 20323 14033
rect 20294 14013 20323 14016
rect 20524 14033 20553 14036
rect 20524 14016 20530 14033
rect 20547 14016 20553 14033
rect 20524 14013 20553 14016
rect 20616 14033 20645 14036
rect 20616 14016 20622 14033
rect 20639 14016 20645 14033
rect 20616 14013 20645 14016
rect 21352 14033 21381 14036
rect 21352 14016 21358 14033
rect 21375 14016 21381 14033
rect 21352 14013 21381 14016
rect 21398 14033 21427 14036
rect 21398 14016 21404 14033
rect 21421 14032 21427 14033
rect 21421 14018 23490 14032
rect 21421 14016 21427 14018
rect 21398 14013 21427 14016
rect 15216 13984 15394 13998
rect 15216 13978 15219 13984
rect 16935 13978 16938 14004
rect 16964 13998 16967 14004
rect 17073 13998 17076 14004
rect 16964 13984 17076 13998
rect 16964 13978 16967 13984
rect 17073 13978 17076 13984
rect 17102 13978 17105 14004
rect 20063 13978 20066 14004
rect 20092 13978 20095 14004
rect 20302 13998 20316 14013
rect 20624 13998 20638 14013
rect 20302 13984 20638 13998
rect 20799 13978 20802 14004
rect 20828 13998 20831 14004
rect 20828 13984 21420 13998
rect 20828 13978 20831 13984
rect 12381 13964 12384 13970
rect 11033 13950 12384 13964
rect 12381 13944 12384 13950
rect 12410 13944 12413 13970
rect 21406 13968 21420 13984
rect 21489 13978 21492 14004
rect 21518 13998 21521 14004
rect 21536 13999 21565 14002
rect 21536 13998 21542 13999
rect 21518 13984 21542 13998
rect 21518 13978 21521 13984
rect 21536 13982 21542 13984
rect 21559 13982 21565 13999
rect 21536 13979 21565 13982
rect 20570 13965 20599 13968
rect 20570 13948 20576 13965
rect 20593 13964 20599 13965
rect 21398 13965 21427 13968
rect 20593 13950 21374 13964
rect 20593 13948 20599 13950
rect 20570 13945 20599 13948
rect 5205 13930 5208 13936
rect 4524 13916 5208 13930
rect 5205 13910 5208 13916
rect 5234 13910 5237 13936
rect 6401 13910 6404 13936
rect 6430 13910 6433 13936
rect 9622 13931 9651 13934
rect 9622 13914 9628 13931
rect 9645 13930 9651 13931
rect 9667 13930 9670 13936
rect 9645 13916 9670 13930
rect 9645 13914 9651 13916
rect 9622 13911 9651 13914
rect 9667 13910 9670 13916
rect 9696 13910 9699 13936
rect 14589 13910 14592 13936
rect 14618 13930 14621 13936
rect 15234 13931 15263 13934
rect 15234 13930 15240 13931
rect 14618 13916 15240 13930
rect 14618 13910 14621 13916
rect 15234 13914 15240 13916
rect 15257 13914 15263 13931
rect 15234 13911 15263 13914
rect 20063 13910 20066 13936
rect 20092 13930 20095 13936
rect 20615 13930 20618 13936
rect 20092 13916 20618 13930
rect 20092 13910 20095 13916
rect 20615 13910 20618 13916
rect 20644 13910 20647 13936
rect 21360 13930 21374 13950
rect 21398 13948 21404 13965
rect 21421 13948 21427 13965
rect 21398 13945 21427 13948
rect 22915 13930 22918 13936
rect 21360 13916 22918 13930
rect 22915 13910 22918 13916
rect 22944 13910 22947 13936
rect 23476 13930 23490 14018
rect 24387 14012 24390 14038
rect 24416 14032 24419 14038
rect 26089 14032 26092 14038
rect 26118 14036 26121 14038
rect 27294 14036 27308 14086
rect 27423 14080 27426 14086
rect 27452 14080 27455 14106
rect 27515 14100 27518 14106
rect 27509 14080 27518 14100
rect 27544 14080 27547 14106
rect 27509 14047 27523 14080
rect 28325 14067 28354 14070
rect 28325 14050 28331 14067
rect 28348 14066 28354 14067
rect 28348 14052 28458 14066
rect 28348 14050 28354 14052
rect 28325 14047 28354 14050
rect 27494 14044 27523 14047
rect 26118 14033 26136 14036
rect 24416 14018 26092 14032
rect 24416 14012 24419 14018
rect 26089 14012 26092 14018
rect 26130 14016 26136 14033
rect 26118 14013 26136 14016
rect 26987 14033 27016 14036
rect 26987 14016 26993 14033
rect 27010 14032 27016 14033
rect 27240 14033 27269 14036
rect 27240 14032 27246 14033
rect 27010 14018 27246 14032
rect 27010 14016 27016 14018
rect 26987 14013 27016 14016
rect 27240 14016 27246 14018
rect 27263 14016 27269 14033
rect 27240 14013 27269 14016
rect 27294 14033 27326 14036
rect 27294 14016 27303 14033
rect 27320 14016 27326 14033
rect 27294 14013 27326 14016
rect 26118 14012 26121 14013
rect 25951 13978 25954 14004
rect 25980 13978 25983 14004
rect 27101 13978 27104 14004
rect 27130 13998 27133 14004
rect 27294 13998 27308 14013
rect 27390 14012 27393 14038
rect 27419 14012 27422 14038
rect 27439 14028 27468 14031
rect 27439 14011 27445 14028
rect 27462 14011 27468 14028
rect 27494 14027 27500 14044
rect 27517 14027 27523 14044
rect 28444 14038 28458 14052
rect 27561 14036 27564 14038
rect 27494 14024 27523 14027
rect 27552 14033 27564 14036
rect 27552 14016 27558 14033
rect 27552 14013 27564 14016
rect 27561 14012 27564 14013
rect 27590 14012 27593 14038
rect 28251 14012 28254 14038
rect 28280 14036 28283 14038
rect 28280 14033 28298 14036
rect 28292 14016 28298 14033
rect 28280 14013 28298 14016
rect 28280 14012 28283 14013
rect 28435 14012 28438 14038
rect 28464 14012 28467 14038
rect 27439 14008 27468 14011
rect 27130 13984 27308 13998
rect 27130 13978 27133 13984
rect 27147 13944 27150 13970
rect 27176 13964 27179 13970
rect 27285 13964 27288 13970
rect 27176 13950 27288 13964
rect 27176 13944 27179 13950
rect 27285 13944 27288 13950
rect 27314 13964 27317 13970
rect 27447 13964 27461 14008
rect 27699 13978 27702 14004
rect 27728 13998 27731 14004
rect 28067 13998 28070 14004
rect 27728 13984 28070 13998
rect 27728 13978 27731 13984
rect 28067 13978 28070 13984
rect 28096 13998 28099 14004
rect 28114 13999 28143 14002
rect 28114 13998 28120 13999
rect 28096 13984 28120 13998
rect 28096 13978 28099 13984
rect 28114 13982 28120 13984
rect 28137 13982 28143 13999
rect 28114 13979 28143 13982
rect 27314 13950 27461 13964
rect 27314 13944 27317 13950
rect 26227 13930 26230 13936
rect 23476 13916 26230 13930
rect 26227 13910 26230 13916
rect 26256 13910 26259 13936
rect 27239 13910 27242 13936
rect 27268 13910 27271 13936
rect 28987 13910 28990 13936
rect 29016 13930 29019 13936
rect 29149 13931 29178 13934
rect 29149 13930 29155 13931
rect 29016 13916 29155 13930
rect 29016 13910 29019 13916
rect 29149 13914 29155 13916
rect 29172 13914 29178 13931
rect 29149 13911 29178 13914
rect 3036 13848 29992 13896
rect 6195 13829 6224 13832
rect 6195 13812 6201 13829
rect 6218 13828 6224 13829
rect 6263 13828 6266 13834
rect 6218 13814 6266 13828
rect 6218 13812 6224 13814
rect 6195 13809 6224 13812
rect 6263 13808 6266 13814
rect 6292 13808 6295 13834
rect 9507 13829 9536 13832
rect 9507 13812 9513 13829
rect 9530 13828 9536 13829
rect 9621 13828 9624 13834
rect 9530 13814 9624 13828
rect 9530 13812 9536 13814
rect 9507 13809 9536 13812
rect 9621 13808 9624 13814
rect 9650 13808 9653 13834
rect 10771 13828 10774 13834
rect 10688 13814 10774 13828
rect 7643 13740 7646 13766
rect 7672 13760 7675 13766
rect 8471 13760 8474 13766
rect 7672 13746 8474 13760
rect 7672 13740 7675 13746
rect 8471 13740 8474 13746
rect 8500 13740 8503 13766
rect 5160 13727 5189 13730
rect 5160 13710 5166 13727
rect 5183 13726 5189 13727
rect 5205 13726 5208 13732
rect 5183 13712 5208 13726
rect 5183 13710 5189 13712
rect 5160 13707 5189 13710
rect 5205 13706 5208 13712
rect 5234 13726 5237 13732
rect 5711 13726 5714 13732
rect 5234 13712 5714 13726
rect 5234 13706 5237 13712
rect 5711 13706 5714 13712
rect 5740 13706 5743 13732
rect 8609 13706 8612 13732
rect 8638 13730 8641 13732
rect 8638 13727 8662 13730
rect 8638 13710 8639 13727
rect 8656 13726 8662 13727
rect 8885 13726 8888 13732
rect 8656 13712 8888 13726
rect 8656 13710 8662 13712
rect 8638 13707 8662 13710
rect 8638 13706 8641 13707
rect 8885 13706 8888 13712
rect 8914 13706 8917 13732
rect 10035 13706 10038 13732
rect 10064 13726 10067 13732
rect 10688 13730 10702 13814
rect 10771 13808 10774 13814
rect 10800 13808 10803 13834
rect 11715 13829 11744 13832
rect 11715 13812 11721 13829
rect 11738 13828 11744 13829
rect 12197 13828 12200 13834
rect 11738 13814 12200 13828
rect 11738 13812 11744 13814
rect 11715 13809 11744 13812
rect 12197 13808 12200 13814
rect 12226 13808 12229 13834
rect 15211 13829 15240 13832
rect 15211 13812 15217 13829
rect 15234 13828 15240 13829
rect 15417 13828 15420 13834
rect 15234 13814 15420 13828
rect 15234 13812 15240 13814
rect 15211 13809 15240 13812
rect 15417 13808 15420 13814
rect 15446 13808 15449 13834
rect 16751 13808 16754 13834
rect 16780 13808 16783 13834
rect 22317 13808 22320 13834
rect 22346 13828 22349 13834
rect 22685 13828 22688 13834
rect 22346 13814 22688 13828
rect 22346 13808 22349 13814
rect 22685 13808 22688 13814
rect 22714 13808 22717 13834
rect 25515 13829 25544 13832
rect 25515 13812 25521 13829
rect 25538 13828 25544 13829
rect 25767 13828 25770 13834
rect 25538 13814 25770 13828
rect 25538 13812 25544 13814
rect 25515 13809 25544 13812
rect 25767 13808 25770 13814
rect 25796 13808 25799 13834
rect 27055 13808 27058 13834
rect 27084 13828 27087 13834
rect 27561 13828 27564 13834
rect 27084 13814 27564 13828
rect 27084 13808 27087 13814
rect 27561 13808 27564 13814
rect 27590 13808 27593 13834
rect 23008 13795 23037 13798
rect 23008 13778 23014 13795
rect 23031 13794 23037 13795
rect 24065 13794 24068 13800
rect 23031 13780 24068 13794
rect 23031 13778 23037 13780
rect 23008 13775 23037 13778
rect 24065 13774 24068 13780
rect 24094 13774 24097 13800
rect 25353 13774 25356 13800
rect 25382 13794 25385 13800
rect 26826 13795 26855 13798
rect 26826 13794 26832 13795
rect 25382 13780 26832 13794
rect 25382 13774 25385 13780
rect 26826 13778 26832 13780
rect 26849 13778 26855 13795
rect 26826 13775 26855 13778
rect 16797 13740 16800 13766
rect 16826 13740 16829 13766
rect 17073 13740 17076 13766
rect 17102 13760 17105 13766
rect 18684 13761 18713 13764
rect 18684 13760 18690 13761
rect 17102 13746 18690 13760
rect 17102 13740 17105 13746
rect 18684 13744 18690 13746
rect 18707 13744 18713 13761
rect 18684 13741 18713 13744
rect 24341 13740 24344 13766
rect 24370 13760 24373 13766
rect 24480 13761 24509 13764
rect 24480 13760 24486 13761
rect 24370 13746 24486 13760
rect 24370 13740 24373 13746
rect 24480 13744 24486 13746
rect 24503 13744 24509 13761
rect 26964 13761 26993 13764
rect 24480 13741 24509 13744
rect 26788 13746 26894 13760
rect 10680 13727 10709 13730
rect 10680 13726 10686 13727
rect 10064 13712 10686 13726
rect 10064 13706 10067 13712
rect 10680 13710 10686 13712
rect 10703 13710 10709 13727
rect 10680 13707 10709 13710
rect 10725 13706 10728 13732
rect 10754 13726 10757 13732
rect 10841 13727 10870 13730
rect 10841 13726 10847 13727
rect 10754 13712 10847 13726
rect 10754 13706 10757 13712
rect 10841 13710 10847 13712
rect 10864 13726 10870 13727
rect 11001 13726 11004 13732
rect 10864 13712 11004 13726
rect 10864 13710 10870 13712
rect 10841 13707 10870 13710
rect 11001 13706 11004 13712
rect 11030 13706 11033 13732
rect 14175 13706 14178 13732
rect 14204 13706 14207 13732
rect 14331 13727 14360 13730
rect 14331 13726 14337 13727
rect 14230 13712 14337 13726
rect 5113 13672 5116 13698
rect 5142 13692 5145 13698
rect 5389 13696 5392 13698
rect 5320 13693 5349 13696
rect 5320 13692 5326 13693
rect 5142 13678 5326 13692
rect 5142 13672 5145 13678
rect 5320 13676 5326 13678
rect 5343 13676 5349 13693
rect 5320 13673 5349 13676
rect 5371 13693 5392 13696
rect 5371 13676 5377 13693
rect 5371 13673 5392 13676
rect 5389 13672 5392 13673
rect 5418 13672 5421 13698
rect 8683 13693 8712 13696
rect 8683 13676 8689 13693
rect 8706 13692 8712 13693
rect 8747 13692 8750 13698
rect 8706 13678 8750 13692
rect 8706 13676 8712 13678
rect 8683 13673 8712 13676
rect 8747 13672 8750 13678
rect 8776 13672 8779 13698
rect 10909 13696 10912 13698
rect 10891 13693 10912 13696
rect 10891 13676 10897 13693
rect 10891 13673 10912 13676
rect 10909 13672 10912 13673
rect 10938 13672 10941 13698
rect 12933 13672 12936 13698
rect 12962 13692 12965 13698
rect 14230 13692 14244 13712
rect 14331 13710 14337 13712
rect 14354 13726 14360 13727
rect 14497 13726 14500 13732
rect 14354 13712 14500 13726
rect 14354 13710 14360 13712
rect 14331 13707 14360 13710
rect 14497 13706 14500 13712
rect 14526 13706 14529 13732
rect 15923 13706 15926 13732
rect 15952 13726 15955 13732
rect 16660 13727 16689 13730
rect 16660 13726 16666 13727
rect 15952 13712 16666 13726
rect 15952 13706 15955 13712
rect 16660 13710 16666 13712
rect 16683 13710 16689 13727
rect 16660 13707 16689 13710
rect 16706 13727 16735 13730
rect 16706 13710 16712 13727
rect 16729 13726 16735 13727
rect 17809 13726 17812 13732
rect 16729 13712 17812 13726
rect 16729 13710 16735 13712
rect 16706 13707 16735 13710
rect 17809 13706 17812 13712
rect 17838 13706 17841 13732
rect 23099 13706 23102 13732
rect 23128 13706 23131 13732
rect 23145 13706 23148 13732
rect 23174 13706 23177 13732
rect 24387 13706 24390 13732
rect 24416 13726 24419 13732
rect 26788 13730 26802 13746
rect 24635 13727 24664 13730
rect 24635 13726 24641 13727
rect 24416 13712 24641 13726
rect 24416 13706 24419 13712
rect 24635 13710 24641 13712
rect 24658 13710 24664 13727
rect 24635 13707 24664 13710
rect 26780 13727 26809 13730
rect 26780 13710 26786 13727
rect 26803 13710 26809 13727
rect 26780 13707 26809 13710
rect 26825 13706 26828 13732
rect 26854 13706 26857 13732
rect 26880 13726 26894 13746
rect 26964 13744 26970 13761
rect 26987 13760 26993 13761
rect 27239 13760 27242 13766
rect 26987 13746 27242 13760
rect 26987 13744 26993 13746
rect 26964 13741 26993 13744
rect 27239 13740 27242 13746
rect 27268 13740 27271 13766
rect 28620 13761 28649 13764
rect 28620 13744 28626 13761
rect 28643 13744 28649 13761
rect 28620 13741 28649 13744
rect 27147 13726 27150 13732
rect 26880 13712 27150 13726
rect 27147 13706 27150 13712
rect 27176 13706 27179 13732
rect 28628 13726 28642 13741
rect 27754 13712 28642 13726
rect 28822 13727 28851 13730
rect 12962 13678 14244 13692
rect 14387 13693 14416 13696
rect 12962 13672 12965 13678
rect 14387 13676 14393 13693
rect 14410 13692 14416 13693
rect 14451 13692 14454 13698
rect 14410 13678 14454 13692
rect 14410 13676 14416 13678
rect 14387 13673 14416 13676
rect 14451 13672 14454 13678
rect 14480 13672 14483 13698
rect 18821 13696 18824 13698
rect 18818 13673 18824 13696
rect 18821 13672 18824 13673
rect 18850 13672 18853 13698
rect 21489 13672 21492 13698
rect 21518 13692 21521 13698
rect 24709 13696 24712 13698
rect 23008 13693 23037 13696
rect 23008 13692 23014 13693
rect 21518 13678 23014 13692
rect 21518 13672 21521 13678
rect 23008 13676 23014 13678
rect 23031 13676 23037 13693
rect 23008 13673 23037 13676
rect 24691 13693 24712 13696
rect 24691 13676 24697 13693
rect 24691 13673 24712 13676
rect 24709 13672 24712 13673
rect 24738 13672 24741 13698
rect 27754 13692 27768 13712
rect 28822 13710 28828 13727
rect 28845 13726 28851 13727
rect 28895 13726 28898 13732
rect 28845 13712 28898 13726
rect 28845 13710 28851 13712
rect 28822 13707 28851 13710
rect 28895 13706 28898 13712
rect 28924 13706 28927 13732
rect 29493 13706 29496 13732
rect 29522 13706 29525 13732
rect 29585 13706 29588 13732
rect 29614 13706 29617 13732
rect 26880 13678 27768 13692
rect 19373 13638 19376 13664
rect 19402 13638 19405 13664
rect 26880 13662 26894 13678
rect 28573 13672 28576 13698
rect 28602 13692 28605 13698
rect 28620 13693 28649 13696
rect 28620 13692 28626 13693
rect 28602 13678 28626 13692
rect 28602 13672 28605 13678
rect 28620 13676 28626 13678
rect 28643 13676 28649 13693
rect 28620 13673 28649 13676
rect 28711 13672 28714 13698
rect 28740 13672 28743 13698
rect 28758 13693 28787 13696
rect 28758 13676 28764 13693
rect 28781 13692 28787 13693
rect 28987 13692 28990 13698
rect 28781 13678 28990 13692
rect 28781 13676 28787 13678
rect 28758 13673 28787 13676
rect 28987 13672 28990 13678
rect 29016 13672 29019 13698
rect 26872 13659 26901 13662
rect 26872 13642 26878 13659
rect 26895 13642 26901 13659
rect 26872 13639 26901 13642
rect 29539 13638 29542 13664
rect 29568 13638 29571 13664
rect 3036 13576 29992 13624
rect 5021 13536 5024 13562
rect 5050 13536 5053 13562
rect 9667 13536 9670 13562
rect 9696 13536 9699 13562
rect 15325 13536 15328 13562
rect 15354 13560 15357 13562
rect 15354 13557 15378 13560
rect 15354 13540 15355 13557
rect 15372 13540 15378 13557
rect 15354 13537 15378 13540
rect 15354 13536 15357 13537
rect 16291 13536 16294 13562
rect 16320 13536 16323 13562
rect 19373 13556 19376 13562
rect 18462 13542 19376 13556
rect 3549 13526 3552 13528
rect 3531 13523 3552 13526
rect 3531 13506 3537 13523
rect 3531 13503 3552 13506
rect 3549 13502 3552 13503
rect 3578 13502 3581 13528
rect 4355 13523 4384 13526
rect 4355 13506 4361 13523
rect 4378 13522 4384 13523
rect 4746 13523 4775 13526
rect 4746 13522 4752 13523
rect 4378 13508 4752 13522
rect 4378 13506 4384 13508
rect 4355 13503 4384 13506
rect 4746 13506 4752 13508
rect 4769 13506 4775 13523
rect 5030 13522 5044 13536
rect 5068 13523 5097 13526
rect 5068 13522 5074 13523
rect 5030 13508 5074 13522
rect 4746 13503 4775 13506
rect 5068 13506 5074 13508
rect 5091 13506 5097 13523
rect 5068 13503 5097 13506
rect 6953 13502 6956 13528
rect 6982 13522 6985 13528
rect 7068 13523 7097 13526
rect 7068 13522 7074 13523
rect 6982 13508 7074 13522
rect 6982 13502 6985 13508
rect 7068 13506 7074 13508
rect 7091 13506 7097 13523
rect 7068 13503 7097 13506
rect 7119 13523 7148 13526
rect 7119 13506 7125 13523
rect 7142 13522 7148 13523
rect 7183 13522 7186 13528
rect 7142 13508 7186 13522
rect 7142 13506 7148 13508
rect 7119 13503 7148 13506
rect 7183 13502 7186 13508
rect 7212 13502 7215 13528
rect 8287 13502 8290 13528
rect 8316 13522 8319 13528
rect 9576 13523 9605 13526
rect 9576 13522 9582 13523
rect 8316 13508 9582 13522
rect 8316 13502 8319 13508
rect 9576 13506 9582 13508
rect 9599 13506 9605 13523
rect 9576 13503 9605 13506
rect 9622 13523 9651 13526
rect 9622 13506 9628 13523
rect 9645 13522 9651 13523
rect 9851 13522 9854 13528
rect 9645 13508 9854 13522
rect 9645 13506 9651 13508
rect 9622 13503 9651 13506
rect 9851 13502 9854 13508
rect 9880 13502 9883 13528
rect 10265 13526 10268 13528
rect 10247 13523 10268 13526
rect 10247 13506 10253 13523
rect 10247 13503 10268 13506
rect 10265 13502 10268 13503
rect 10294 13502 10297 13528
rect 11645 13502 11648 13528
rect 11674 13522 11677 13528
rect 14543 13526 14546 13528
rect 13007 13523 13036 13526
rect 13007 13522 13013 13523
rect 11674 13508 13013 13522
rect 11674 13502 11677 13508
rect 13007 13506 13013 13508
rect 13030 13522 13036 13523
rect 14525 13523 14546 13526
rect 13030 13506 13048 13522
rect 13007 13503 13048 13506
rect 14525 13506 14531 13523
rect 14525 13503 14546 13506
rect 3319 13468 3322 13494
rect 3348 13468 3351 13494
rect 3457 13468 3460 13494
rect 3486 13492 3489 13494
rect 3486 13489 3504 13492
rect 3498 13472 3504 13489
rect 3486 13469 3504 13472
rect 3486 13468 3489 13469
rect 4607 13468 4610 13494
rect 4636 13468 4639 13494
rect 4700 13489 4729 13492
rect 4700 13472 4706 13489
rect 4723 13472 4729 13489
rect 4700 13469 4729 13472
rect 4810 13489 4839 13492
rect 4810 13472 4816 13489
rect 4833 13488 4839 13489
rect 5021 13488 5024 13494
rect 4833 13474 5024 13488
rect 4833 13472 4839 13474
rect 4810 13469 4839 13472
rect 4708 13420 4722 13469
rect 5021 13468 5024 13474
rect 5050 13468 5053 13494
rect 5159 13468 5162 13494
rect 5188 13468 5191 13494
rect 5206 13489 5235 13492
rect 5206 13472 5212 13489
rect 5229 13472 5235 13489
rect 5206 13469 5235 13472
rect 4746 13455 4775 13458
rect 4746 13438 4752 13455
rect 4769 13454 4775 13455
rect 5214 13454 5228 13469
rect 6309 13468 6312 13494
rect 6338 13488 6341 13494
rect 9162 13489 9191 13492
rect 9162 13488 9168 13489
rect 6338 13474 9168 13488
rect 6338 13468 6341 13474
rect 9162 13472 9168 13474
rect 9185 13472 9191 13489
rect 9162 13469 9191 13472
rect 4769 13440 5228 13454
rect 4769 13438 4775 13440
rect 4746 13435 4775 13438
rect 6861 13434 6864 13460
rect 6890 13454 6893 13460
rect 6908 13455 6937 13458
rect 6908 13454 6914 13455
rect 6890 13440 6914 13454
rect 6890 13434 6893 13440
rect 6908 13438 6914 13440
rect 6931 13438 6937 13455
rect 9170 13454 9184 13469
rect 9253 13468 9256 13494
rect 9282 13468 9285 13494
rect 10197 13489 10226 13492
rect 10197 13472 10203 13489
rect 10220 13488 10226 13489
rect 10311 13488 10314 13494
rect 10220 13474 10314 13488
rect 10220 13472 10226 13474
rect 10197 13469 10226 13472
rect 10311 13468 10314 13474
rect 10340 13488 10343 13494
rect 10725 13488 10728 13494
rect 10340 13474 10728 13488
rect 10340 13468 10343 13474
rect 10725 13468 10728 13474
rect 10754 13468 10757 13494
rect 12336 13489 12365 13492
rect 12336 13488 12342 13489
rect 11033 13474 12342 13488
rect 9170 13440 9552 13454
rect 6908 13435 6937 13438
rect 5113 13420 5116 13426
rect 4708 13406 5116 13420
rect 5113 13400 5116 13406
rect 5142 13420 5145 13426
rect 8103 13420 8106 13426
rect 5142 13406 6930 13420
rect 5142 13400 5145 13406
rect 5206 13387 5235 13390
rect 5206 13370 5212 13387
rect 5229 13386 5235 13387
rect 6171 13386 6174 13392
rect 5229 13372 6174 13386
rect 5229 13370 5235 13372
rect 5206 13367 5235 13370
rect 6171 13366 6174 13372
rect 6200 13366 6203 13392
rect 6916 13386 6930 13406
rect 7721 13406 8106 13420
rect 7721 13386 7735 13406
rect 8103 13400 8106 13406
rect 8132 13400 8135 13426
rect 9208 13421 9237 13424
rect 9208 13404 9214 13421
rect 9231 13420 9237 13421
rect 9484 13421 9513 13424
rect 9484 13420 9490 13421
rect 9231 13406 9490 13420
rect 9231 13404 9237 13406
rect 9208 13401 9237 13404
rect 9484 13404 9490 13406
rect 9507 13404 9513 13421
rect 9538 13420 9552 13440
rect 10035 13434 10038 13460
rect 10064 13434 10067 13460
rect 9538 13406 10058 13420
rect 9484 13401 9513 13404
rect 6916 13372 7735 13386
rect 7943 13387 7972 13390
rect 7943 13370 7949 13387
rect 7966 13386 7972 13387
rect 8011 13386 8014 13392
rect 7966 13372 8014 13386
rect 7966 13370 7972 13372
rect 7943 13367 7972 13370
rect 8011 13366 8014 13372
rect 8040 13366 8043 13392
rect 9760 13387 9789 13390
rect 9760 13370 9766 13387
rect 9783 13386 9789 13387
rect 9943 13386 9946 13392
rect 9783 13372 9946 13386
rect 9783 13370 9789 13372
rect 9760 13367 9789 13370
rect 9943 13366 9946 13372
rect 9972 13366 9975 13392
rect 10044 13386 10058 13406
rect 11033 13386 11047 13474
rect 12336 13472 12342 13474
rect 12359 13472 12365 13489
rect 12336 13469 12365 13472
rect 12344 13454 12358 13469
rect 12427 13468 12430 13494
rect 12456 13468 12459 13494
rect 12519 13468 12522 13494
rect 12548 13488 12551 13494
rect 12933 13488 12936 13494
rect 12962 13492 12965 13494
rect 12962 13489 12980 13492
rect 12548 13474 12936 13488
rect 12548 13468 12551 13474
rect 12933 13468 12936 13474
rect 12974 13472 12980 13489
rect 13034 13488 13048 13503
rect 14543 13502 14546 13503
rect 14572 13502 14575 13528
rect 17073 13522 17076 13528
rect 15610 13508 17076 13522
rect 14359 13488 14362 13494
rect 13034 13474 14362 13488
rect 12962 13469 12980 13472
rect 12962 13468 12965 13469
rect 14359 13468 14362 13474
rect 14388 13468 14391 13494
rect 14451 13468 14454 13494
rect 14480 13492 14483 13494
rect 14480 13489 14498 13492
rect 14492 13472 14498 13489
rect 14480 13469 14498 13472
rect 14480 13468 14483 13469
rect 15610 13460 15624 13508
rect 17073 13502 17076 13508
rect 17102 13502 17105 13528
rect 17717 13502 17720 13528
rect 17746 13522 17749 13528
rect 17855 13522 17858 13528
rect 17746 13508 17858 13522
rect 17746 13502 17749 13508
rect 17855 13502 17858 13508
rect 17884 13522 17887 13528
rect 18462 13522 18476 13542
rect 19373 13536 19376 13542
rect 19402 13536 19405 13562
rect 27033 13557 27062 13560
rect 27033 13540 27039 13557
rect 27056 13556 27062 13557
rect 27423 13556 27426 13562
rect 27056 13542 27426 13556
rect 27056 13540 27062 13542
rect 27033 13537 27062 13540
rect 27423 13536 27426 13542
rect 27452 13536 27455 13562
rect 19511 13522 19514 13528
rect 17884 13508 18476 13522
rect 17884 13502 17887 13508
rect 15736 13489 15765 13492
rect 15736 13472 15742 13489
rect 15759 13488 15765 13489
rect 16015 13488 16018 13494
rect 15759 13474 16018 13488
rect 15759 13472 15765 13474
rect 15736 13469 15765 13472
rect 16015 13468 16018 13474
rect 16044 13468 16047 13494
rect 18315 13468 18318 13494
rect 18344 13488 18347 13494
rect 18462 13492 18476 13508
rect 18876 13508 19514 13522
rect 18408 13489 18437 13492
rect 18408 13488 18414 13489
rect 18344 13474 18414 13488
rect 18344 13468 18347 13474
rect 18408 13472 18414 13474
rect 18431 13472 18437 13489
rect 18408 13469 18437 13472
rect 18455 13489 18484 13492
rect 18455 13472 18461 13489
rect 18478 13472 18484 13489
rect 18455 13469 18484 13472
rect 18826 13489 18855 13492
rect 18826 13472 18832 13489
rect 18849 13483 18855 13489
rect 18876 13483 18890 13508
rect 19511 13502 19514 13508
rect 19540 13502 19543 13528
rect 26209 13523 26238 13526
rect 26209 13506 26215 13523
rect 26232 13522 26238 13523
rect 26232 13508 26342 13522
rect 26232 13506 26238 13508
rect 26209 13503 26238 13506
rect 26328 13494 26342 13508
rect 18849 13472 18890 13483
rect 18826 13469 18890 13472
rect 19051 13468 19054 13494
rect 19080 13468 19083 13494
rect 24204 13489 24233 13492
rect 24204 13472 24210 13489
rect 24227 13488 24233 13489
rect 25353 13488 25356 13494
rect 24227 13474 25356 13488
rect 24227 13472 24233 13474
rect 24204 13469 24233 13472
rect 25353 13468 25356 13474
rect 25382 13468 25385 13494
rect 25997 13468 26000 13494
rect 26026 13468 26029 13494
rect 26135 13468 26138 13494
rect 26164 13492 26167 13494
rect 26164 13489 26182 13492
rect 26176 13472 26182 13489
rect 26164 13469 26182 13472
rect 26164 13468 26167 13469
rect 26319 13468 26322 13494
rect 26348 13488 26351 13494
rect 27009 13488 27012 13494
rect 26348 13474 27012 13488
rect 26348 13468 26351 13474
rect 27009 13468 27012 13474
rect 27038 13468 27041 13494
rect 12749 13454 12752 13460
rect 12344 13440 12752 13454
rect 12749 13434 12752 13440
rect 12778 13434 12781 13460
rect 12795 13434 12798 13460
rect 12824 13434 12827 13460
rect 14175 13434 14178 13460
rect 14204 13454 14207 13460
rect 14313 13454 14316 13460
rect 14204 13440 14316 13454
rect 14204 13434 14207 13440
rect 14313 13434 14316 13440
rect 14342 13434 14345 13460
rect 15601 13434 15604 13460
rect 15630 13434 15633 13460
rect 18960 13455 18989 13458
rect 18960 13438 18966 13455
rect 18983 13454 18989 13455
rect 20063 13454 20066 13460
rect 18983 13440 20066 13454
rect 18983 13438 18989 13440
rect 18960 13435 18989 13438
rect 20063 13434 20066 13440
rect 20092 13434 20095 13460
rect 21397 13434 21400 13460
rect 21426 13454 21429 13460
rect 21581 13454 21584 13460
rect 21426 13440 21584 13454
rect 21426 13434 21429 13440
rect 21581 13434 21584 13440
rect 21610 13434 21613 13460
rect 24157 13434 24160 13460
rect 24186 13434 24189 13460
rect 24296 13455 24325 13458
rect 24296 13438 24302 13455
rect 24319 13438 24325 13455
rect 24296 13435 24325 13438
rect 18592 13421 18621 13424
rect 18592 13404 18598 13421
rect 18615 13420 18621 13421
rect 18729 13420 18732 13426
rect 18615 13406 18732 13420
rect 18615 13404 18621 13406
rect 18592 13401 18621 13404
rect 18729 13400 18732 13406
rect 18758 13400 18761 13426
rect 18775 13400 18778 13426
rect 18804 13420 18807 13426
rect 19006 13421 19035 13424
rect 19006 13420 19012 13421
rect 18804 13406 19012 13420
rect 18804 13400 18807 13406
rect 19006 13404 19012 13406
rect 19029 13404 19035 13421
rect 19006 13401 19035 13404
rect 21351 13400 21354 13426
rect 21380 13420 21383 13426
rect 24304 13420 24318 13435
rect 21380 13406 24318 13420
rect 21380 13400 21383 13406
rect 10044 13372 11047 13386
rect 11071 13387 11100 13390
rect 11071 13370 11077 13387
rect 11094 13386 11100 13387
rect 11875 13386 11878 13392
rect 11094 13372 11878 13386
rect 11094 13370 11100 13372
rect 11071 13367 11100 13370
rect 11875 13366 11878 13372
rect 11904 13366 11907 13392
rect 12382 13387 12411 13390
rect 12382 13370 12388 13387
rect 12405 13386 12411 13387
rect 12473 13386 12476 13392
rect 12405 13372 12476 13386
rect 12405 13370 12411 13372
rect 12382 13367 12411 13370
rect 12473 13366 12476 13372
rect 12502 13366 12505 13392
rect 13831 13387 13860 13390
rect 13831 13370 13837 13387
rect 13854 13386 13860 13387
rect 14681 13386 14684 13392
rect 13854 13372 14684 13386
rect 13854 13370 13860 13372
rect 13831 13367 13860 13370
rect 14681 13366 14684 13372
rect 14710 13366 14713 13392
rect 16521 13366 16524 13392
rect 16550 13386 16553 13392
rect 18891 13387 18920 13390
rect 18891 13386 18897 13387
rect 16550 13372 18897 13386
rect 16550 13366 16553 13372
rect 18891 13370 18897 13372
rect 18914 13370 18920 13387
rect 18891 13367 18920 13370
rect 24249 13366 24252 13392
rect 24278 13366 24281 13392
rect 3036 13304 29992 13352
rect 3319 13284 3322 13290
rect 3144 13270 3322 13284
rect 3144 13222 3158 13270
rect 3319 13264 3322 13270
rect 3348 13264 3351 13290
rect 4171 13285 4200 13288
rect 4171 13268 4177 13285
rect 4194 13284 4200 13285
rect 4607 13284 4610 13290
rect 4194 13270 4610 13284
rect 4194 13268 4200 13270
rect 4171 13265 4200 13268
rect 4607 13264 4610 13270
rect 4636 13264 4639 13290
rect 4837 13264 4840 13290
rect 4866 13284 4869 13290
rect 8195 13284 8198 13290
rect 4866 13270 8198 13284
rect 4866 13264 4869 13270
rect 8195 13264 8198 13270
rect 8224 13264 8227 13290
rect 10081 13264 10084 13290
rect 10110 13284 10113 13290
rect 10110 13270 12404 13284
rect 10110 13264 10113 13270
rect 7874 13251 7903 13254
rect 7874 13234 7880 13251
rect 7897 13250 7903 13251
rect 8287 13250 8290 13256
rect 7897 13236 8290 13250
rect 7897 13234 7903 13236
rect 7874 13231 7903 13234
rect 8287 13230 8290 13236
rect 8316 13230 8319 13256
rect 3135 13196 3138 13222
rect 3164 13196 3167 13222
rect 4792 13217 4821 13220
rect 4792 13200 4798 13217
rect 4815 13216 4821 13217
rect 5159 13216 5162 13222
rect 4815 13202 5162 13216
rect 4815 13200 4821 13202
rect 4792 13197 4821 13200
rect 5159 13196 5162 13202
rect 5188 13196 5191 13222
rect 5205 13196 5208 13222
rect 5234 13216 5237 13222
rect 5343 13216 5346 13222
rect 5234 13202 5346 13216
rect 5234 13196 5237 13202
rect 5343 13196 5346 13202
rect 5372 13196 5375 13222
rect 6203 13202 8724 13216
rect 3297 13183 3326 13186
rect 3297 13166 3303 13183
rect 3320 13182 3326 13183
rect 3457 13182 3460 13188
rect 3320 13168 3460 13182
rect 3320 13166 3326 13168
rect 3297 13163 3326 13166
rect 3457 13162 3460 13168
rect 3486 13162 3489 13188
rect 4745 13162 4748 13188
rect 4774 13162 4777 13188
rect 4837 13162 4840 13188
rect 4866 13186 4869 13188
rect 4866 13182 4870 13186
rect 4866 13168 4888 13182
rect 4866 13163 4870 13168
rect 4866 13162 4869 13163
rect 5389 13162 5392 13188
rect 5418 13182 5421 13188
rect 6203 13182 6217 13202
rect 5418 13168 6217 13182
rect 5418 13162 5421 13168
rect 3365 13152 3368 13154
rect 3347 13149 3368 13152
rect 3347 13132 3353 13149
rect 3347 13129 3368 13132
rect 3365 13128 3368 13129
rect 3394 13128 3397 13154
rect 4653 13128 4656 13154
rect 4682 13128 4685 13154
rect 4791 13128 4794 13154
rect 4820 13128 4823 13154
rect 5297 13128 5300 13154
rect 5326 13148 5329 13154
rect 5505 13149 5534 13152
rect 5505 13148 5511 13149
rect 5326 13134 5511 13148
rect 5326 13128 5329 13134
rect 5505 13132 5511 13134
rect 5528 13132 5534 13149
rect 5505 13129 5534 13132
rect 5555 13149 5584 13152
rect 5555 13132 5561 13149
rect 5578 13148 5584 13149
rect 5674 13148 5688 13168
rect 7873 13162 7876 13188
rect 7902 13162 7905 13188
rect 7919 13162 7922 13188
rect 7948 13186 7951 13188
rect 7948 13183 7960 13186
rect 7954 13166 7960 13183
rect 7948 13163 7960 13166
rect 7948 13162 7951 13163
rect 8011 13162 8014 13188
rect 8040 13184 8043 13188
rect 8040 13181 8054 13184
rect 8048 13164 8054 13181
rect 8040 13162 8054 13164
rect 8086 13162 8089 13188
rect 8115 13162 8118 13188
rect 8195 13186 8198 13188
rect 8186 13183 8198 13186
rect 8135 13173 8164 13176
rect 8025 13161 8054 13162
rect 8135 13156 8141 13173
rect 8158 13156 8164 13173
rect 8186 13166 8192 13183
rect 8186 13163 8198 13166
rect 8195 13162 8198 13163
rect 8224 13162 8227 13188
rect 8471 13162 8474 13188
rect 8500 13182 8503 13188
rect 8656 13183 8685 13186
rect 8656 13182 8662 13183
rect 8500 13168 8662 13182
rect 8500 13162 8503 13168
rect 8656 13166 8662 13168
rect 8679 13166 8685 13183
rect 8710 13182 8724 13202
rect 10035 13196 10038 13222
rect 10064 13216 10067 13222
rect 11416 13217 11445 13220
rect 11416 13216 11422 13217
rect 10064 13202 11422 13216
rect 10064 13196 10067 13202
rect 11416 13200 11422 13202
rect 11439 13200 11445 13217
rect 12390 13216 12404 13270
rect 12427 13264 12430 13290
rect 12456 13288 12459 13290
rect 12456 13285 12480 13288
rect 12456 13268 12457 13285
rect 12474 13268 12480 13285
rect 12456 13265 12480 13268
rect 12456 13264 12459 13265
rect 12749 13264 12752 13290
rect 12778 13284 12781 13290
rect 15877 13284 15880 13290
rect 12778 13270 15880 13284
rect 12778 13264 12781 13270
rect 14681 13230 14684 13256
rect 14710 13230 14713 13256
rect 12390 13202 13324 13216
rect 11416 13197 11445 13200
rect 11047 13182 11050 13188
rect 8710 13168 11050 13182
rect 8656 13163 8685 13166
rect 8135 13153 8164 13156
rect 5578 13134 5688 13148
rect 5578 13132 5584 13134
rect 5555 13129 5584 13132
rect 8143 13120 8157 13153
rect 8609 13128 8612 13154
rect 8638 13148 8641 13154
rect 8894 13152 8908 13168
rect 11047 13162 11050 13168
rect 11076 13162 11079 13188
rect 11571 13183 11600 13186
rect 11571 13182 11577 13183
rect 11102 13168 11577 13182
rect 8816 13149 8845 13152
rect 8816 13148 8822 13149
rect 8638 13134 8822 13148
rect 8638 13128 8641 13134
rect 8816 13132 8822 13134
rect 8839 13132 8845 13149
rect 8816 13129 8845 13132
rect 8867 13149 8908 13152
rect 8867 13132 8873 13149
rect 8890 13134 8908 13149
rect 8890 13132 8896 13134
rect 8867 13129 8896 13132
rect 11001 13128 11004 13154
rect 11030 13148 11033 13154
rect 11102 13148 11116 13168
rect 11571 13166 11577 13168
rect 11594 13166 11600 13183
rect 11571 13163 11600 13166
rect 12795 13162 12798 13188
rect 12824 13182 12827 13188
rect 13256 13183 13285 13186
rect 13256 13182 13262 13183
rect 12824 13168 13262 13182
rect 12824 13162 12827 13168
rect 13256 13166 13262 13168
rect 13279 13166 13285 13183
rect 13310 13182 13324 13202
rect 13577 13182 13580 13188
rect 13310 13168 13580 13182
rect 13256 13163 13285 13166
rect 13577 13162 13580 13168
rect 13606 13162 13609 13188
rect 14497 13162 14500 13188
rect 14526 13182 14529 13188
rect 14635 13186 14638 13188
rect 14544 13183 14573 13186
rect 14544 13182 14550 13183
rect 14526 13168 14550 13182
rect 14526 13162 14529 13168
rect 14544 13166 14550 13168
rect 14567 13166 14573 13183
rect 14544 13163 14573 13166
rect 14621 13183 14638 13186
rect 14621 13166 14627 13183
rect 14621 13163 14638 13166
rect 14635 13162 14638 13163
rect 14664 13162 14667 13188
rect 14690 13184 14704 13230
rect 14751 13192 14765 13270
rect 15877 13264 15880 13270
rect 15906 13264 15909 13290
rect 16015 13264 16018 13290
rect 16044 13284 16047 13290
rect 16062 13285 16091 13288
rect 16062 13284 16068 13285
rect 16044 13270 16068 13284
rect 16044 13264 16047 13270
rect 16062 13268 16068 13270
rect 16085 13268 16091 13285
rect 16062 13265 16091 13268
rect 18776 13285 18805 13288
rect 18776 13268 18782 13285
rect 18799 13284 18805 13285
rect 18821 13284 18824 13290
rect 18799 13270 18824 13284
rect 18799 13268 18805 13270
rect 18776 13265 18805 13268
rect 18821 13264 18824 13270
rect 18850 13264 18853 13290
rect 24157 13264 24160 13290
rect 24186 13284 24189 13290
rect 29539 13284 29542 13290
rect 24186 13270 29542 13284
rect 24186 13264 24189 13270
rect 29539 13264 29542 13270
rect 29568 13264 29571 13290
rect 14819 13230 14822 13256
rect 14848 13230 14851 13256
rect 16338 13251 16367 13254
rect 16338 13250 16344 13251
rect 15978 13236 16344 13250
rect 14828 13192 14842 13230
rect 15978 13220 15992 13236
rect 16338 13234 16344 13236
rect 16361 13234 16367 13251
rect 16338 13231 16367 13234
rect 23145 13230 23148 13256
rect 23174 13250 23177 13256
rect 28757 13250 28760 13256
rect 23174 13236 28760 13250
rect 23174 13230 23177 13236
rect 28757 13230 28760 13236
rect 28786 13230 28789 13256
rect 15970 13217 15999 13220
rect 15970 13200 15976 13217
rect 15993 13200 15999 13217
rect 15970 13197 15999 13200
rect 16108 13217 16137 13220
rect 16108 13200 16114 13217
rect 16131 13216 16137 13217
rect 16935 13216 16938 13222
rect 16131 13202 16938 13216
rect 16131 13200 16137 13202
rect 16108 13197 16137 13200
rect 16935 13196 16938 13202
rect 16964 13216 16967 13222
rect 16964 13202 18798 13216
rect 16964 13196 16967 13202
rect 14743 13189 14772 13192
rect 14690 13181 14724 13184
rect 14690 13165 14701 13181
rect 14695 13164 14701 13165
rect 14718 13164 14724 13181
rect 14743 13172 14749 13189
rect 14766 13172 14772 13189
rect 14743 13169 14772 13172
rect 14805 13189 14842 13192
rect 14805 13172 14811 13189
rect 14828 13173 14842 13189
rect 14856 13183 14885 13186
rect 14828 13172 14834 13173
rect 14805 13169 14834 13172
rect 11030 13134 11116 13148
rect 11030 13128 11033 13134
rect 11277 13128 11280 13154
rect 11306 13148 11309 13154
rect 11645 13152 11648 13154
rect 11627 13149 11648 13152
rect 11627 13148 11633 13149
rect 11306 13134 11633 13148
rect 11306 13128 11309 13134
rect 11627 13132 11633 13134
rect 11627 13129 11648 13132
rect 11645 13128 11648 13129
rect 11674 13128 11677 13154
rect 12933 13128 12936 13154
rect 12962 13148 12965 13154
rect 13416 13149 13445 13152
rect 13416 13148 13422 13149
rect 12962 13134 13422 13148
rect 12962 13128 12965 13134
rect 13416 13132 13422 13134
rect 13439 13132 13445 13149
rect 13416 13129 13445 13132
rect 13467 13149 13496 13152
rect 13467 13132 13473 13149
rect 13490 13148 13496 13149
rect 13586 13148 13600 13162
rect 14695 13161 14724 13164
rect 14856 13166 14862 13183
rect 14879 13182 14885 13183
rect 14957 13182 14960 13188
rect 14879 13168 14960 13182
rect 14879 13166 14885 13168
rect 14856 13163 14885 13166
rect 14957 13162 14960 13168
rect 14986 13162 14989 13188
rect 16016 13183 16045 13186
rect 16016 13166 16022 13183
rect 16039 13166 16045 13183
rect 16016 13163 16045 13166
rect 16024 13148 16038 13163
rect 16291 13162 16294 13188
rect 16320 13182 16323 13188
rect 16338 13183 16367 13186
rect 16338 13182 16344 13183
rect 16320 13168 16344 13182
rect 16320 13162 16323 13168
rect 16338 13166 16344 13168
rect 16361 13166 16367 13183
rect 16338 13163 16367 13166
rect 16476 13183 16505 13186
rect 16476 13166 16482 13183
rect 16499 13182 16505 13183
rect 16567 13182 16570 13188
rect 16499 13168 16570 13182
rect 16499 13166 16505 13168
rect 16476 13163 16505 13166
rect 16567 13162 16570 13168
rect 16596 13162 16599 13188
rect 18638 13183 18667 13186
rect 18638 13166 18644 13183
rect 18661 13182 18667 13183
rect 18683 13182 18686 13188
rect 18661 13168 18686 13182
rect 18661 13166 18667 13168
rect 18638 13163 18667 13166
rect 18683 13162 18686 13168
rect 18712 13162 18715 13188
rect 18729 13162 18732 13188
rect 18758 13162 18761 13188
rect 18784 13186 18798 13202
rect 20845 13196 20848 13222
rect 20874 13216 20877 13222
rect 20874 13202 21282 13216
rect 20874 13196 20877 13202
rect 18776 13183 18805 13186
rect 18776 13166 18782 13183
rect 18799 13166 18805 13183
rect 18776 13163 18805 13166
rect 21213 13162 21216 13188
rect 21242 13162 21245 13188
rect 21268 13182 21282 13202
rect 21375 13183 21404 13186
rect 21375 13182 21381 13183
rect 21268 13168 21381 13182
rect 21375 13166 21381 13168
rect 21398 13166 21404 13183
rect 21375 13163 21404 13166
rect 21535 13162 21538 13188
rect 21564 13162 21567 13188
rect 21903 13162 21906 13188
rect 21932 13182 21935 13188
rect 22823 13182 22826 13188
rect 21932 13168 22826 13182
rect 21932 13162 21935 13168
rect 22823 13162 22826 13168
rect 22852 13162 22855 13188
rect 19281 13148 19284 13154
rect 13490 13134 13600 13148
rect 14483 13134 14612 13148
rect 16024 13134 19284 13148
rect 13490 13132 13496 13134
rect 13467 13129 13496 13132
rect 6355 13094 6358 13120
rect 6384 13118 6387 13120
rect 6384 13115 6408 13118
rect 6384 13098 6385 13115
rect 6402 13098 6408 13115
rect 8143 13100 8152 13120
rect 6384 13095 6408 13098
rect 6384 13094 6387 13095
rect 8149 13094 8152 13100
rect 8178 13094 8181 13120
rect 9691 13115 9720 13118
rect 9691 13098 9697 13115
rect 9714 13114 9720 13115
rect 9759 13114 9762 13120
rect 9714 13100 9762 13114
rect 9714 13098 9720 13100
rect 9691 13095 9720 13098
rect 9759 13094 9762 13100
rect 9788 13094 9791 13120
rect 14291 13115 14320 13118
rect 14291 13098 14297 13115
rect 14314 13114 14320 13115
rect 14483 13114 14497 13134
rect 14314 13100 14497 13114
rect 14314 13098 14320 13100
rect 14291 13095 14320 13098
rect 14543 13094 14546 13120
rect 14572 13094 14575 13120
rect 14598 13114 14612 13134
rect 19281 13128 19284 13134
rect 19310 13128 19313 13154
rect 21425 13149 21454 13152
rect 21425 13132 21431 13149
rect 21448 13148 21454 13149
rect 21544 13148 21558 13162
rect 21448 13134 21558 13148
rect 21448 13132 21454 13134
rect 21425 13129 21454 13132
rect 14819 13114 14822 13120
rect 14598 13100 14822 13114
rect 14819 13094 14822 13100
rect 14848 13094 14851 13120
rect 16430 13115 16459 13118
rect 16430 13098 16436 13115
rect 16453 13114 16459 13115
rect 17165 13114 17168 13120
rect 16453 13100 17168 13114
rect 16453 13098 16459 13100
rect 16430 13095 16459 13098
rect 17165 13094 17168 13100
rect 17194 13094 17197 13120
rect 22249 13115 22278 13118
rect 22249 13098 22255 13115
rect 22272 13114 22278 13115
rect 22869 13114 22872 13120
rect 22272 13100 22872 13114
rect 22272 13098 22278 13100
rect 22249 13095 22278 13098
rect 22869 13094 22872 13100
rect 22898 13094 22901 13120
rect 3036 13032 29992 13080
rect 4677 13013 4706 13016
rect 4677 12996 4683 13013
rect 4700 13012 4706 13013
rect 4791 13012 4794 13018
rect 4700 12998 4794 13012
rect 4700 12996 4706 12998
rect 4677 12993 4706 12996
rect 4791 12992 4794 12998
rect 4820 12992 4823 13018
rect 5297 12992 5300 13018
rect 5326 13012 5329 13018
rect 5619 13012 5622 13018
rect 5326 12998 5622 13012
rect 5326 12992 5329 12998
rect 5619 12992 5622 12998
rect 5648 12992 5651 13018
rect 7989 13013 8018 13016
rect 7989 12996 7995 13013
rect 8012 13012 8018 13013
rect 8149 13012 8152 13018
rect 8012 12998 8152 13012
rect 8012 12996 8018 12998
rect 7989 12993 8018 12996
rect 8149 12992 8152 12998
rect 8178 12992 8181 13018
rect 11968 13013 11997 13016
rect 11968 12996 11974 13013
rect 11991 13012 11997 13013
rect 12336 13013 12365 13016
rect 12336 13012 12342 13013
rect 11991 12998 12342 13012
rect 11991 12996 11997 12998
rect 11968 12993 11997 12996
rect 12336 12996 12342 12998
rect 12359 12996 12365 13013
rect 12336 12993 12365 12996
rect 12381 12992 12384 13018
rect 12410 12992 12413 13018
rect 13831 13013 13860 13016
rect 13831 12996 13837 13013
rect 13854 13012 13860 13013
rect 14497 13012 14500 13018
rect 13854 12998 14500 13012
rect 13854 12996 13860 12998
rect 13831 12993 13860 12996
rect 14497 12992 14500 12998
rect 14526 12992 14529 13018
rect 19281 12992 19284 13018
rect 19310 13012 19313 13018
rect 19328 13013 19357 13016
rect 19328 13012 19334 13013
rect 19310 12998 19334 13012
rect 19310 12992 19313 12998
rect 19328 12996 19334 12998
rect 19351 12996 19357 13013
rect 19328 12993 19357 12996
rect 22777 12992 22780 13018
rect 22806 13012 22809 13018
rect 22806 12998 22938 13012
rect 22806 12992 22809 12998
rect 3871 12982 3874 12984
rect 3853 12979 3874 12982
rect 3853 12962 3859 12979
rect 3900 12978 3903 12984
rect 3900 12964 3986 12978
rect 3853 12959 3874 12962
rect 3871 12958 3874 12959
rect 3900 12958 3903 12964
rect 3457 12924 3460 12950
rect 3486 12944 3489 12950
rect 3803 12945 3832 12948
rect 3803 12944 3809 12945
rect 3486 12930 3809 12944
rect 3486 12924 3489 12930
rect 3803 12928 3809 12930
rect 3826 12944 3832 12945
rect 3917 12944 3920 12950
rect 3826 12930 3920 12944
rect 3826 12928 3832 12930
rect 3803 12925 3832 12928
rect 3917 12924 3920 12930
rect 3946 12924 3949 12950
rect 3972 12944 3986 12964
rect 6309 12958 6312 12984
rect 6338 12958 6341 12984
rect 6355 12958 6358 12984
rect 6384 12958 6387 12984
rect 6447 12978 6450 12984
rect 6410 12964 6450 12978
rect 3972 12930 5826 12944
rect 3135 12890 3138 12916
rect 3164 12910 3167 12916
rect 3642 12911 3671 12914
rect 3642 12910 3648 12911
rect 3164 12896 3648 12910
rect 3164 12890 3167 12896
rect 3642 12894 3648 12896
rect 3665 12894 3671 12911
rect 3642 12891 3671 12894
rect 5812 12876 5826 12930
rect 6171 12924 6174 12950
rect 6200 12924 6203 12950
rect 6217 12924 6220 12950
rect 6246 12924 6249 12950
rect 6410 12948 6424 12964
rect 6447 12958 6450 12964
rect 6476 12958 6479 12984
rect 7165 12979 7194 12982
rect 7165 12978 7171 12979
rect 6916 12964 7171 12978
rect 6402 12945 6431 12948
rect 6402 12928 6408 12945
rect 6425 12928 6431 12945
rect 6402 12925 6431 12928
rect 6448 12911 6477 12914
rect 6448 12894 6454 12911
rect 6471 12910 6477 12911
rect 6493 12910 6496 12916
rect 6471 12896 6496 12910
rect 6471 12894 6477 12896
rect 6448 12891 6477 12894
rect 6493 12890 6496 12896
rect 6522 12890 6525 12916
rect 6916 12876 6930 12964
rect 7165 12962 7171 12964
rect 7188 12978 7194 12979
rect 7188 12964 7298 12978
rect 7188 12962 7194 12964
rect 7165 12959 7194 12962
rect 7091 12924 7094 12950
rect 7120 12948 7123 12950
rect 7120 12945 7138 12948
rect 7132 12928 7138 12945
rect 7284 12944 7298 12964
rect 10081 12958 10084 12984
rect 10110 12978 10113 12984
rect 13025 12982 13028 12984
rect 10243 12979 10272 12982
rect 10243 12978 10249 12979
rect 10110 12964 10249 12978
rect 10110 12958 10113 12964
rect 10243 12962 10249 12964
rect 10266 12962 10272 12979
rect 10243 12959 10272 12962
rect 11071 12979 11100 12982
rect 11071 12962 11077 12979
rect 11094 12978 11100 12979
rect 13007 12979 13028 12982
rect 11094 12964 11806 12978
rect 11094 12962 11100 12964
rect 11071 12959 11100 12962
rect 9115 12944 9118 12950
rect 7284 12930 9118 12944
rect 7120 12925 7138 12928
rect 7120 12924 7123 12925
rect 9115 12924 9118 12930
rect 9144 12924 9147 12950
rect 10197 12945 10226 12948
rect 10197 12928 10203 12945
rect 10220 12944 10226 12945
rect 10311 12944 10314 12950
rect 10220 12930 10314 12944
rect 10220 12928 10226 12930
rect 10197 12925 10226 12928
rect 10311 12924 10314 12930
rect 10340 12924 10343 12950
rect 11737 12924 11740 12950
rect 11766 12924 11769 12950
rect 11792 12948 11806 12964
rect 13007 12962 13013 12979
rect 13007 12959 13028 12962
rect 13025 12958 13028 12959
rect 13054 12958 13057 12984
rect 16429 12978 16432 12984
rect 16162 12964 16432 12978
rect 11792 12945 11824 12948
rect 11792 12930 11801 12945
rect 11795 12928 11801 12930
rect 11818 12928 11824 12945
rect 11795 12925 11824 12928
rect 11875 12924 11878 12950
rect 11904 12948 11907 12950
rect 12059 12948 12062 12950
rect 11904 12945 11918 12948
rect 11912 12928 11918 12945
rect 12050 12945 12062 12948
rect 11904 12925 11918 12928
rect 11951 12940 11980 12943
rect 11904 12924 11907 12925
rect 11951 12923 11957 12940
rect 11974 12923 11980 12940
rect 11951 12920 11980 12923
rect 11999 12940 12028 12943
rect 11999 12923 12005 12940
rect 12022 12938 12028 12940
rect 12022 12923 12036 12938
rect 12050 12928 12056 12945
rect 12050 12925 12062 12928
rect 12059 12924 12062 12925
rect 12088 12924 12091 12950
rect 12243 12924 12246 12950
rect 12272 12944 12275 12950
rect 12290 12945 12319 12948
rect 12290 12944 12296 12945
rect 12272 12930 12296 12944
rect 12272 12924 12275 12930
rect 12290 12928 12296 12930
rect 12313 12928 12319 12945
rect 12290 12925 12319 12928
rect 12473 12924 12476 12950
rect 12502 12924 12505 12950
rect 12933 12924 12936 12950
rect 12962 12948 12965 12950
rect 16162 12948 16176 12964
rect 16429 12958 16432 12964
rect 16458 12978 16461 12984
rect 17441 12978 17444 12984
rect 16458 12964 17444 12978
rect 16458 12958 16461 12964
rect 17441 12958 17444 12964
rect 17470 12958 17473 12984
rect 19235 12958 19238 12984
rect 19264 12958 19267 12984
rect 20799 12978 20802 12984
rect 19336 12964 20802 12978
rect 12962 12945 12980 12948
rect 12974 12928 12980 12945
rect 12962 12925 12980 12928
rect 16154 12945 16183 12948
rect 16154 12928 16160 12945
rect 16177 12928 16183 12945
rect 16154 12925 16183 12928
rect 12962 12924 12965 12925
rect 16475 12924 16478 12950
rect 16504 12924 16507 12950
rect 19190 12945 19219 12948
rect 19190 12928 19196 12945
rect 19213 12944 19219 12945
rect 19336 12944 19350 12964
rect 20799 12958 20802 12964
rect 20828 12958 20831 12984
rect 20845 12958 20848 12984
rect 20874 12978 20877 12984
rect 21029 12982 21032 12984
rect 20960 12979 20989 12982
rect 20960 12978 20966 12979
rect 20874 12964 20966 12978
rect 20874 12958 20877 12964
rect 20960 12962 20966 12964
rect 20983 12962 20989 12979
rect 20960 12959 20989 12962
rect 21011 12979 21032 12982
rect 21011 12962 21017 12979
rect 21011 12959 21032 12962
rect 21029 12958 21032 12959
rect 21058 12958 21061 12984
rect 22823 12978 22826 12984
rect 22815 12958 22826 12978
rect 22852 12958 22855 12984
rect 19213 12930 19350 12944
rect 19213 12928 19219 12930
rect 19190 12925 19219 12928
rect 19373 12924 19376 12950
rect 19402 12924 19405 12950
rect 21835 12945 21864 12948
rect 21835 12928 21841 12945
rect 21858 12944 21864 12945
rect 22594 12945 22623 12948
rect 22594 12944 22600 12945
rect 21858 12930 22600 12944
rect 21858 12928 21864 12930
rect 21835 12925 21864 12928
rect 22594 12928 22600 12930
rect 22617 12928 22623 12945
rect 22594 12925 22623 12928
rect 22639 12924 22642 12950
rect 22668 12948 22671 12950
rect 22745 12948 22774 12951
rect 22668 12945 22680 12948
rect 22745 12946 22751 12948
rect 22674 12928 22680 12945
rect 22668 12925 22680 12928
rect 22696 12932 22751 12946
rect 22668 12924 22671 12925
rect 11999 12920 12036 12923
rect 6954 12911 6983 12914
rect 6954 12894 6960 12911
rect 6977 12894 6983 12911
rect 6954 12891 6983 12894
rect 5812 12862 6930 12876
rect 6861 12822 6864 12848
rect 6890 12842 6893 12848
rect 6962 12842 6976 12891
rect 10035 12890 10038 12916
rect 10064 12890 10067 12916
rect 6890 12828 6976 12842
rect 6890 12822 6893 12828
rect 9023 12822 9026 12848
rect 9052 12842 9055 12848
rect 10265 12842 10268 12848
rect 9052 12828 10268 12842
rect 9052 12822 9055 12828
rect 10265 12822 10268 12828
rect 10294 12822 10297 12848
rect 11959 12842 11973 12920
rect 12022 12876 12036 12920
rect 12795 12890 12798 12916
rect 12824 12890 12827 12916
rect 16522 12911 16551 12914
rect 16522 12894 16528 12911
rect 16545 12910 16551 12911
rect 16567 12910 16570 12916
rect 16545 12896 16570 12910
rect 16545 12894 16551 12896
rect 16522 12891 16551 12894
rect 16567 12890 16570 12896
rect 16596 12910 16599 12916
rect 17073 12910 17076 12916
rect 16596 12896 17076 12910
rect 16596 12890 16599 12896
rect 17073 12890 17076 12896
rect 17102 12890 17105 12916
rect 19281 12890 19284 12916
rect 19310 12890 19313 12916
rect 20800 12911 20829 12914
rect 20800 12894 20806 12911
rect 20823 12894 20829 12911
rect 20800 12891 20829 12894
rect 12059 12876 12062 12882
rect 12022 12862 12062 12876
rect 12059 12856 12062 12862
rect 12088 12856 12091 12882
rect 12390 12862 12818 12876
rect 12390 12842 12404 12862
rect 11959 12828 12404 12842
rect 12427 12822 12430 12848
rect 12456 12822 12459 12848
rect 12804 12842 12818 12862
rect 14819 12842 14822 12848
rect 12804 12828 14822 12842
rect 14819 12822 14822 12828
rect 14848 12822 14851 12848
rect 20808 12842 20822 12891
rect 22271 12890 22274 12916
rect 22300 12910 22303 12916
rect 22696 12910 22710 12932
rect 22745 12931 22751 12932
rect 22768 12931 22774 12948
rect 22815 12943 22829 12958
rect 22924 12950 22938 12998
rect 29493 12992 29496 13018
rect 29522 12992 29525 13018
rect 25859 12958 25862 12984
rect 25888 12978 25891 12984
rect 26067 12979 26096 12982
rect 26067 12978 26073 12979
rect 25888 12964 26073 12978
rect 25888 12958 25891 12964
rect 26067 12962 26073 12964
rect 26090 12962 26096 12979
rect 26067 12959 26096 12962
rect 28113 12958 28116 12984
rect 28142 12978 28145 12984
rect 28251 12978 28254 12984
rect 28142 12964 28254 12978
rect 28142 12958 28145 12964
rect 28251 12958 28254 12964
rect 28280 12978 28283 12984
rect 28366 12979 28395 12982
rect 28366 12978 28372 12979
rect 28280 12964 28372 12978
rect 28280 12958 28283 12964
rect 28366 12962 28372 12964
rect 28389 12962 28395 12979
rect 28366 12959 28395 12962
rect 28417 12979 28446 12982
rect 28417 12962 28423 12979
rect 28440 12978 28446 12979
rect 28440 12964 28550 12978
rect 28440 12962 28446 12964
rect 28417 12959 28446 12962
rect 28536 12950 28550 12964
rect 22915 12948 22918 12950
rect 22906 12945 22918 12948
rect 22745 12928 22774 12931
rect 22807 12940 22836 12943
rect 22807 12923 22813 12940
rect 22830 12923 22836 12940
rect 22807 12920 22836 12923
rect 22855 12940 22884 12943
rect 22855 12923 22861 12940
rect 22878 12938 22884 12940
rect 22878 12923 22892 12938
rect 22906 12928 22912 12945
rect 22906 12925 22918 12928
rect 22915 12924 22918 12925
rect 22944 12924 22947 12950
rect 25629 12924 25632 12950
rect 25658 12944 25661 12950
rect 26021 12945 26050 12948
rect 26021 12944 26027 12945
rect 25658 12930 26027 12944
rect 25658 12924 25661 12930
rect 26021 12928 26027 12930
rect 26044 12944 26050 12945
rect 26135 12944 26138 12950
rect 26044 12930 26138 12944
rect 26044 12928 26050 12930
rect 26021 12925 26050 12928
rect 26135 12924 26138 12930
rect 26164 12924 26167 12950
rect 28527 12924 28530 12950
rect 28556 12924 28559 12950
rect 29401 12924 29404 12950
rect 29430 12944 29433 12950
rect 29494 12945 29523 12948
rect 29494 12944 29500 12945
rect 29430 12930 29500 12944
rect 29430 12924 29433 12930
rect 29494 12928 29500 12930
rect 29517 12928 29523 12945
rect 29494 12925 29523 12928
rect 29539 12924 29542 12950
rect 29568 12948 29571 12950
rect 29568 12945 29580 12948
rect 29574 12928 29580 12945
rect 29568 12925 29580 12928
rect 29568 12924 29571 12925
rect 29631 12924 29634 12950
rect 29660 12948 29663 12950
rect 29660 12945 29684 12948
rect 29660 12928 29661 12945
rect 29678 12928 29684 12945
rect 29660 12925 29684 12928
rect 29660 12924 29663 12925
rect 29706 12924 29709 12950
rect 29735 12924 29738 12950
rect 29815 12948 29818 12950
rect 29755 12945 29784 12948
rect 29755 12928 29761 12945
rect 29778 12928 29784 12945
rect 29755 12925 29784 12928
rect 29806 12945 29818 12948
rect 29806 12928 29812 12945
rect 29806 12925 29818 12928
rect 22855 12920 22892 12923
rect 22300 12896 22710 12910
rect 22300 12890 22303 12896
rect 22878 12882 22892 12920
rect 25860 12911 25889 12914
rect 25860 12894 25866 12911
rect 25883 12894 25889 12911
rect 25860 12891 25889 12894
rect 22869 12856 22872 12882
rect 22898 12856 22901 12882
rect 21213 12842 21216 12848
rect 20808 12828 21216 12842
rect 21213 12822 21216 12828
rect 21242 12822 21245 12848
rect 22593 12822 22596 12848
rect 22622 12822 22625 12848
rect 25537 12822 25540 12848
rect 25566 12842 25569 12848
rect 25868 12842 25882 12891
rect 27837 12890 27840 12916
rect 27866 12910 27869 12916
rect 28067 12910 28070 12916
rect 27866 12896 28070 12910
rect 27866 12890 27869 12896
rect 28067 12890 28070 12896
rect 28096 12910 28099 12916
rect 28206 12911 28235 12914
rect 28206 12910 28212 12911
rect 28096 12896 28212 12910
rect 28096 12890 28099 12896
rect 28206 12894 28212 12896
rect 28229 12894 28235 12911
rect 28206 12891 28235 12894
rect 29241 12911 29270 12914
rect 29241 12894 29247 12911
rect 29264 12910 29270 12911
rect 29763 12910 29777 12925
rect 29815 12924 29818 12925
rect 29844 12924 29847 12950
rect 29264 12896 29777 12910
rect 29264 12894 29270 12896
rect 29241 12891 29270 12894
rect 25997 12842 26000 12848
rect 25566 12828 26000 12842
rect 25566 12822 25569 12828
rect 25997 12822 26000 12828
rect 26026 12822 26029 12848
rect 26895 12843 26924 12846
rect 26895 12826 26901 12843
rect 26918 12842 26924 12843
rect 27331 12842 27334 12848
rect 26918 12828 27334 12842
rect 26918 12826 26924 12828
rect 26895 12823 26924 12826
rect 27331 12822 27334 12828
rect 27360 12822 27363 12848
rect 3036 12760 29992 12808
rect 4171 12741 4200 12744
rect 4171 12724 4177 12741
rect 4194 12740 4200 12741
rect 4653 12740 4656 12746
rect 4194 12726 4656 12740
rect 4194 12724 4200 12726
rect 4171 12721 4200 12724
rect 4653 12720 4656 12726
rect 4682 12720 4685 12746
rect 5343 12740 5346 12746
rect 5214 12726 5346 12740
rect 3135 12652 3138 12678
rect 3164 12652 3167 12678
rect 5214 12676 5228 12726
rect 5343 12720 5346 12726
rect 5372 12720 5375 12746
rect 6217 12720 6220 12746
rect 6246 12744 6249 12746
rect 6246 12741 6270 12744
rect 6246 12724 6247 12741
rect 6264 12724 6270 12741
rect 8333 12740 8336 12746
rect 6246 12721 6270 12724
rect 6456 12726 8336 12740
rect 6246 12720 6249 12721
rect 5206 12673 5235 12676
rect 5206 12656 5212 12673
rect 5229 12656 5235 12673
rect 5206 12653 5235 12656
rect 3297 12639 3326 12642
rect 3297 12622 3303 12639
rect 3320 12638 3326 12639
rect 3457 12638 3460 12644
rect 3320 12624 3460 12638
rect 3320 12622 3326 12624
rect 3297 12619 3326 12622
rect 3457 12618 3460 12624
rect 3486 12618 3489 12644
rect 5251 12618 5254 12644
rect 5280 12638 5283 12644
rect 5405 12639 5434 12642
rect 5405 12638 5411 12639
rect 5280 12624 5411 12638
rect 5280 12618 5283 12624
rect 5405 12622 5411 12624
rect 5428 12638 5434 12639
rect 6456 12638 6470 12726
rect 8333 12720 8336 12726
rect 8362 12740 8365 12746
rect 9139 12741 9168 12744
rect 8362 12726 9092 12740
rect 8362 12720 8365 12726
rect 9078 12706 9092 12726
rect 9139 12724 9145 12741
rect 9162 12740 9168 12741
rect 9253 12740 9256 12746
rect 9162 12726 9256 12740
rect 9162 12724 9168 12726
rect 9139 12721 9168 12724
rect 9253 12720 9256 12726
rect 9282 12720 9285 12746
rect 11277 12740 11280 12746
rect 9653 12726 11280 12740
rect 9653 12706 9667 12726
rect 11277 12720 11280 12726
rect 11306 12720 11309 12746
rect 11899 12741 11928 12744
rect 11899 12724 11905 12741
rect 11922 12740 11928 12741
rect 12059 12740 12062 12746
rect 11922 12726 12062 12740
rect 11922 12724 11928 12726
rect 11899 12721 11928 12724
rect 12059 12720 12062 12726
rect 12088 12720 12091 12746
rect 13992 12741 14021 12744
rect 13992 12724 13998 12741
rect 14015 12740 14021 12741
rect 14037 12740 14040 12746
rect 14015 12726 14040 12740
rect 14015 12724 14021 12726
rect 13992 12721 14021 12724
rect 14037 12720 14040 12726
rect 14066 12720 14069 12746
rect 22271 12744 22274 12746
rect 22249 12741 22274 12744
rect 22249 12724 22255 12741
rect 22272 12724 22274 12741
rect 22249 12721 22274 12724
rect 22271 12720 22274 12721
rect 22300 12720 22303 12746
rect 28873 12741 28902 12744
rect 28873 12724 28879 12741
rect 28896 12740 28902 12741
rect 29539 12740 29542 12746
rect 28896 12726 29542 12740
rect 28896 12724 28902 12726
rect 28873 12721 28902 12724
rect 29539 12720 29542 12726
rect 29568 12720 29571 12746
rect 9078 12692 9667 12706
rect 6861 12652 6864 12678
rect 6890 12672 6893 12678
rect 8104 12673 8133 12676
rect 8104 12672 8110 12673
rect 6890 12658 8110 12672
rect 6890 12652 6893 12658
rect 8104 12656 8110 12658
rect 8127 12656 8133 12673
rect 8104 12653 8133 12656
rect 10035 12652 10038 12678
rect 10064 12672 10067 12678
rect 10864 12673 10893 12676
rect 10864 12672 10870 12673
rect 10064 12658 10870 12672
rect 10064 12652 10067 12658
rect 10864 12656 10870 12658
rect 10887 12656 10893 12673
rect 14589 12672 14592 12678
rect 10864 12653 10893 12656
rect 14506 12658 14592 12672
rect 5428 12624 6470 12638
rect 5428 12622 5434 12624
rect 5405 12619 5434 12622
rect 6493 12618 6496 12644
rect 6522 12618 6525 12644
rect 6632 12639 6661 12642
rect 6632 12622 6638 12639
rect 6655 12638 6661 12639
rect 7229 12638 7232 12644
rect 6655 12624 7232 12638
rect 6655 12622 6661 12624
rect 6632 12619 6661 12622
rect 7229 12618 7232 12624
rect 7258 12618 7261 12644
rect 10311 12618 10314 12644
rect 10340 12638 10343 12644
rect 10449 12638 10452 12644
rect 10340 12624 10452 12638
rect 10340 12618 10343 12624
rect 10449 12618 10452 12624
rect 10478 12638 10481 12644
rect 11019 12639 11048 12642
rect 11019 12638 11025 12639
rect 10478 12624 11025 12638
rect 10478 12618 10481 12624
rect 11019 12622 11025 12624
rect 11042 12622 11048 12639
rect 13025 12638 13028 12644
rect 11019 12619 11048 12622
rect 11194 12624 13028 12638
rect 3347 12605 3376 12608
rect 3347 12588 3353 12605
rect 3370 12604 3376 12605
rect 3411 12604 3414 12610
rect 3370 12590 3414 12604
rect 3370 12588 3376 12590
rect 3347 12585 3376 12588
rect 3411 12584 3414 12590
rect 3440 12584 3443 12610
rect 4745 12584 4748 12610
rect 4774 12604 4777 12610
rect 4975 12604 4978 12610
rect 4774 12590 4978 12604
rect 4774 12584 4777 12590
rect 4975 12584 4978 12590
rect 5004 12584 5007 12610
rect 5366 12605 5395 12608
rect 5366 12604 5372 12605
rect 5260 12590 5372 12604
rect 5260 12576 5274 12590
rect 5366 12588 5372 12590
rect 5389 12588 5395 12605
rect 5366 12585 5395 12588
rect 6586 12605 6615 12608
rect 6586 12588 6592 12605
rect 6609 12604 6615 12605
rect 7413 12604 7416 12610
rect 6609 12590 7416 12604
rect 6609 12588 6615 12590
rect 6586 12585 6615 12588
rect 7413 12584 7416 12590
rect 7442 12584 7445 12610
rect 8149 12584 8152 12610
rect 8178 12604 8181 12610
rect 8333 12608 8336 12610
rect 8264 12605 8293 12608
rect 8264 12604 8270 12605
rect 8178 12590 8270 12604
rect 8178 12584 8181 12590
rect 8264 12588 8270 12590
rect 8287 12588 8293 12605
rect 8264 12585 8293 12588
rect 8315 12605 8336 12608
rect 8315 12588 8321 12605
rect 8315 12585 8336 12588
rect 8333 12584 8336 12585
rect 8362 12584 8365 12610
rect 9115 12584 9118 12610
rect 9144 12604 9147 12610
rect 11075 12605 11104 12608
rect 11075 12604 11081 12605
rect 9144 12590 11081 12604
rect 9144 12584 9147 12590
rect 11075 12588 11081 12590
rect 11098 12604 11104 12605
rect 11194 12604 11208 12624
rect 13025 12618 13028 12624
rect 13054 12618 13057 12644
rect 14506 12642 14520 12658
rect 14589 12652 14592 12658
rect 14618 12652 14621 12678
rect 16567 12672 16570 12678
rect 15863 12658 16570 12672
rect 14498 12639 14527 12642
rect 14498 12622 14504 12639
rect 14521 12622 14527 12639
rect 14498 12619 14527 12622
rect 14543 12618 14546 12644
rect 14572 12618 14575 12644
rect 14681 12618 14684 12644
rect 14710 12618 14713 12644
rect 15693 12618 15696 12644
rect 15722 12618 15725 12644
rect 15786 12639 15815 12642
rect 15786 12622 15792 12639
rect 15809 12638 15815 12639
rect 15863 12638 15877 12658
rect 16567 12652 16570 12658
rect 16596 12652 16599 12678
rect 19879 12652 19882 12678
rect 19908 12672 19911 12678
rect 19908 12658 20316 12672
rect 19908 12652 19911 12658
rect 15809 12624 15877 12638
rect 15809 12622 15815 12624
rect 15786 12619 15815 12622
rect 16429 12618 16432 12644
rect 16458 12618 16461 12644
rect 16521 12618 16524 12644
rect 16550 12618 16553 12644
rect 16752 12639 16781 12642
rect 16752 12622 16758 12639
rect 16775 12622 16781 12639
rect 16752 12619 16781 12622
rect 11098 12590 11208 12604
rect 11098 12588 11104 12590
rect 11075 12585 11104 12588
rect 13899 12584 13902 12610
rect 13928 12584 13931 12610
rect 16291 12584 16294 12610
rect 16320 12604 16323 12610
rect 16475 12604 16478 12610
rect 16320 12590 16478 12604
rect 16320 12584 16323 12590
rect 16475 12584 16478 12590
rect 16504 12604 16507 12610
rect 16760 12604 16774 12619
rect 19511 12618 19514 12644
rect 19540 12638 19543 12644
rect 19971 12638 19974 12644
rect 19540 12624 19974 12638
rect 19540 12618 19543 12624
rect 19971 12618 19974 12624
rect 20000 12638 20003 12644
rect 20302 12642 20316 12658
rect 21213 12652 21216 12678
rect 21242 12652 21245 12678
rect 22409 12652 22412 12678
rect 22438 12672 22441 12678
rect 22639 12672 22642 12678
rect 22438 12658 22642 12672
rect 22438 12652 22441 12658
rect 22639 12652 22642 12658
rect 22668 12652 22671 12678
rect 25583 12652 25586 12678
rect 25612 12672 25615 12678
rect 26273 12672 26276 12678
rect 25612 12658 26276 12672
rect 25612 12652 25615 12658
rect 26273 12652 26276 12658
rect 26302 12652 26305 12678
rect 20064 12639 20093 12642
rect 20064 12638 20070 12639
rect 20000 12624 20070 12638
rect 20000 12618 20003 12624
rect 20064 12622 20070 12624
rect 20087 12622 20093 12639
rect 20064 12619 20093 12622
rect 20294 12639 20323 12642
rect 20294 12622 20300 12639
rect 20317 12622 20323 12639
rect 20845 12638 20848 12644
rect 20294 12619 20323 12622
rect 20693 12624 20848 12638
rect 16504 12590 16774 12604
rect 16504 12584 16507 12590
rect 20431 12584 20434 12610
rect 20460 12584 20463 12610
rect 20477 12584 20480 12610
rect 20506 12604 20509 12610
rect 20693 12604 20707 12624
rect 20845 12618 20848 12624
rect 20874 12638 20877 12644
rect 21369 12639 21398 12642
rect 21369 12638 21375 12639
rect 20874 12624 21375 12638
rect 20874 12618 20877 12624
rect 21369 12622 21375 12624
rect 21392 12622 21398 12639
rect 21369 12619 21398 12622
rect 21413 12639 21442 12642
rect 21413 12622 21419 12639
rect 21436 12638 21442 12639
rect 21627 12638 21630 12644
rect 21436 12624 21630 12638
rect 21436 12622 21442 12624
rect 21413 12619 21442 12622
rect 21627 12618 21630 12624
rect 21656 12618 21659 12644
rect 27837 12618 27840 12644
rect 27866 12618 27869 12644
rect 27999 12639 28028 12642
rect 27999 12622 28005 12639
rect 28022 12638 28028 12639
rect 28113 12638 28116 12644
rect 28022 12624 28116 12638
rect 28022 12622 28028 12624
rect 27999 12619 28028 12622
rect 28113 12618 28116 12624
rect 28142 12618 28145 12644
rect 28159 12618 28162 12644
rect 28188 12618 28191 12644
rect 28067 12608 28070 12610
rect 20506 12590 20707 12604
rect 28049 12605 28070 12608
rect 20506 12584 20509 12590
rect 28049 12588 28055 12605
rect 28096 12604 28099 12610
rect 28168 12604 28182 12618
rect 28096 12590 28182 12604
rect 28049 12585 28070 12588
rect 28067 12584 28070 12585
rect 28096 12584 28099 12590
rect 3917 12550 3920 12576
rect 3946 12570 3949 12576
rect 5251 12570 5254 12576
rect 3946 12556 5254 12570
rect 3946 12550 3949 12556
rect 5251 12550 5254 12556
rect 5280 12550 5283 12576
rect 6539 12550 6542 12576
rect 6568 12550 6571 12576
rect 11691 12550 11694 12576
rect 11720 12570 11723 12576
rect 12611 12570 12614 12576
rect 11720 12556 12614 12570
rect 11720 12550 11723 12556
rect 12611 12550 12614 12556
rect 12640 12550 12643 12576
rect 13991 12550 13994 12576
rect 14020 12574 14023 12576
rect 14020 12571 14029 12574
rect 14023 12554 14029 12571
rect 14020 12551 14029 12554
rect 14084 12571 14113 12574
rect 14084 12554 14090 12571
rect 14107 12570 14113 12571
rect 14590 12571 14619 12574
rect 14590 12570 14596 12571
rect 14107 12556 14596 12570
rect 14107 12554 14113 12556
rect 14084 12551 14113 12554
rect 14590 12554 14596 12556
rect 14613 12554 14619 12571
rect 14590 12551 14619 12554
rect 14682 12571 14711 12574
rect 14682 12554 14688 12571
rect 14705 12570 14711 12571
rect 14727 12570 14730 12576
rect 14705 12556 14730 12570
rect 14705 12554 14711 12556
rect 14682 12551 14711 12554
rect 14020 12550 14023 12551
rect 14727 12550 14730 12556
rect 14756 12550 14759 12576
rect 15739 12550 15742 12576
rect 15768 12550 15771 12576
rect 17165 12550 17168 12576
rect 17194 12570 17197 12576
rect 18315 12570 18318 12576
rect 17194 12556 18318 12570
rect 17194 12550 17197 12556
rect 18315 12550 18318 12556
rect 18344 12550 18347 12576
rect 28297 12550 28300 12576
rect 28326 12570 28329 12576
rect 28389 12570 28392 12576
rect 28326 12556 28392 12570
rect 28326 12550 28329 12556
rect 28389 12550 28392 12556
rect 28418 12550 28421 12576
rect 3036 12488 29992 12536
rect 5251 12448 5254 12474
rect 5280 12468 5283 12474
rect 5619 12468 5622 12474
rect 5280 12454 5622 12468
rect 5280 12448 5283 12454
rect 5619 12448 5622 12454
rect 5648 12468 5651 12474
rect 5941 12468 5944 12474
rect 5648 12454 5944 12468
rect 5648 12448 5651 12454
rect 5941 12448 5944 12454
rect 5970 12448 5973 12474
rect 10403 12448 10406 12474
rect 10432 12468 10435 12474
rect 11691 12468 11694 12474
rect 10432 12454 11694 12468
rect 10432 12448 10435 12454
rect 11691 12448 11694 12454
rect 11720 12448 11723 12474
rect 12114 12469 12143 12472
rect 12114 12468 12120 12469
rect 11746 12454 12120 12468
rect 3135 12414 3138 12440
rect 3164 12434 3167 12440
rect 4745 12438 4748 12440
rect 4727 12435 4748 12438
rect 3164 12420 4170 12434
rect 3164 12414 3167 12420
rect 4156 12366 4170 12420
rect 4727 12418 4733 12435
rect 4727 12415 4748 12418
rect 4745 12414 4748 12415
rect 4774 12414 4777 12440
rect 6907 12414 6910 12440
rect 6936 12434 6939 12440
rect 7069 12435 7098 12438
rect 7069 12434 7075 12435
rect 6936 12420 7075 12434
rect 6936 12414 6939 12420
rect 7069 12418 7075 12420
rect 7092 12418 7098 12435
rect 7069 12415 7098 12418
rect 8149 12414 8152 12440
rect 8178 12434 8181 12440
rect 8609 12434 8612 12440
rect 8178 12420 8612 12434
rect 8178 12414 8181 12420
rect 8609 12414 8612 12420
rect 8638 12434 8641 12440
rect 9023 12438 9026 12440
rect 8954 12435 8983 12438
rect 8954 12434 8960 12435
rect 8638 12420 8960 12434
rect 8638 12414 8641 12420
rect 8954 12418 8960 12420
rect 8977 12418 8983 12435
rect 8954 12415 8983 12418
rect 9005 12435 9026 12438
rect 9005 12418 9011 12435
rect 9005 12415 9026 12418
rect 9023 12414 9026 12415
rect 9052 12414 9055 12440
rect 11746 12434 11760 12454
rect 12114 12452 12120 12454
rect 12137 12452 12143 12469
rect 12114 12449 12143 12452
rect 12198 12469 12227 12472
rect 12198 12452 12204 12469
rect 12221 12468 12227 12469
rect 12381 12468 12384 12474
rect 12221 12454 12384 12468
rect 12221 12452 12227 12454
rect 12198 12449 12227 12452
rect 12381 12448 12384 12454
rect 12410 12448 12413 12474
rect 14819 12448 14822 12474
rect 14848 12468 14851 12474
rect 16337 12468 16340 12474
rect 14848 12454 16340 12468
rect 14848 12448 14851 12454
rect 16337 12448 16340 12454
rect 16366 12448 16369 12474
rect 23974 12469 24003 12472
rect 17818 12454 18430 12468
rect 11608 12420 11760 12434
rect 4677 12401 4706 12404
rect 4677 12384 4683 12401
rect 4700 12400 4706 12401
rect 6539 12400 6542 12406
rect 4700 12386 6542 12400
rect 4700 12384 4706 12386
rect 4677 12381 4706 12384
rect 6539 12380 6542 12386
rect 6568 12380 6571 12406
rect 6861 12380 6864 12406
rect 6890 12380 6893 12406
rect 7023 12401 7052 12404
rect 7023 12384 7029 12401
rect 7046 12400 7052 12401
rect 7137 12400 7140 12406
rect 7046 12386 7140 12400
rect 7046 12384 7052 12386
rect 7023 12381 7052 12384
rect 7137 12380 7140 12386
rect 7166 12380 7169 12406
rect 7873 12380 7876 12406
rect 7902 12404 7905 12406
rect 7902 12401 7926 12404
rect 7902 12384 7903 12401
rect 7920 12384 7926 12401
rect 7902 12381 7926 12384
rect 7902 12380 7905 12381
rect 8471 12380 8474 12406
rect 8500 12400 8503 12406
rect 8794 12401 8823 12404
rect 8794 12400 8800 12401
rect 8500 12386 8800 12400
rect 8500 12380 8503 12386
rect 8794 12384 8800 12386
rect 8817 12400 8823 12401
rect 10035 12400 10038 12406
rect 8817 12386 10038 12400
rect 8817 12384 8823 12386
rect 8794 12381 8823 12384
rect 10035 12380 10038 12386
rect 10064 12400 10067 12406
rect 10082 12401 10111 12404
rect 10082 12400 10088 12401
rect 10064 12386 10088 12400
rect 10064 12380 10067 12386
rect 10082 12384 10088 12386
rect 10105 12384 10111 12401
rect 10082 12381 10111 12384
rect 11553 12380 11556 12406
rect 11582 12380 11585 12406
rect 4515 12366 4518 12372
rect 4156 12352 4518 12366
rect 4515 12346 4518 12352
rect 4544 12346 4547 12372
rect 10863 12346 10866 12372
rect 10892 12346 10895 12372
rect 11608 12370 11622 12420
rect 12013 12414 12016 12440
rect 12042 12414 12045 12440
rect 12611 12414 12614 12440
rect 12640 12434 12643 12440
rect 12773 12435 12802 12438
rect 12773 12434 12779 12435
rect 12640 12420 12779 12434
rect 12640 12414 12643 12420
rect 12773 12418 12779 12420
rect 12796 12418 12802 12435
rect 14474 12435 14503 12438
rect 14474 12434 14480 12435
rect 12773 12415 12802 12418
rect 13586 12420 14480 12434
rect 11645 12380 11648 12406
rect 11674 12380 11677 12406
rect 11691 12380 11694 12406
rect 11720 12380 11723 12406
rect 11737 12380 11740 12406
rect 11766 12404 11769 12406
rect 11766 12400 11770 12404
rect 12727 12401 12756 12404
rect 11766 12386 11788 12400
rect 11766 12381 11770 12386
rect 12727 12384 12733 12401
rect 12750 12400 12756 12401
rect 12887 12400 12890 12406
rect 12750 12386 12890 12400
rect 12750 12384 12756 12386
rect 12727 12381 12756 12384
rect 11766 12380 11769 12381
rect 12887 12380 12890 12386
rect 12916 12400 12919 12406
rect 13586 12400 13600 12420
rect 14474 12418 14480 12420
rect 14497 12418 14503 12435
rect 14474 12415 14503 12418
rect 14525 12435 14554 12438
rect 14525 12418 14531 12435
rect 14548 12434 14554 12435
rect 14589 12434 14592 12440
rect 14548 12420 14592 12434
rect 14548 12418 14554 12420
rect 14525 12415 14554 12418
rect 14589 12414 14592 12420
rect 14618 12414 14621 12440
rect 15739 12438 15742 12440
rect 15736 12434 15742 12438
rect 15719 12420 15742 12434
rect 15736 12415 15742 12420
rect 15739 12414 15742 12415
rect 15768 12414 15771 12440
rect 17073 12414 17076 12440
rect 17102 12434 17105 12440
rect 17102 12420 17326 12434
rect 17102 12414 17105 12420
rect 15601 12400 15604 12406
rect 12916 12386 13600 12400
rect 14322 12386 15604 12400
rect 12916 12380 12919 12386
rect 14322 12372 14336 12386
rect 15601 12380 15604 12386
rect 15630 12380 15633 12406
rect 17027 12380 17030 12406
rect 17056 12400 17059 12406
rect 17165 12400 17168 12406
rect 17056 12386 17168 12400
rect 17056 12380 17059 12386
rect 17165 12380 17168 12386
rect 17194 12380 17197 12406
rect 17211 12380 17214 12406
rect 17240 12380 17243 12406
rect 17261 12396 17290 12399
rect 17261 12379 17267 12396
rect 17284 12379 17290 12396
rect 17261 12376 17290 12379
rect 11600 12367 11629 12370
rect 11600 12350 11606 12367
rect 11623 12350 11629 12367
rect 11600 12347 11629 12350
rect 12566 12367 12595 12370
rect 12566 12350 12572 12367
rect 12589 12350 12595 12367
rect 12566 12347 12595 12350
rect 5435 12278 5438 12304
rect 5464 12298 5467 12304
rect 5551 12299 5580 12302
rect 5551 12298 5557 12299
rect 5464 12284 5557 12298
rect 5464 12278 5467 12284
rect 5551 12282 5557 12284
rect 5574 12282 5580 12299
rect 5551 12279 5580 12282
rect 8931 12278 8934 12304
rect 8960 12298 8963 12304
rect 9829 12299 9858 12302
rect 9829 12298 9835 12299
rect 8960 12284 9835 12298
rect 8960 12278 8963 12284
rect 9829 12282 9835 12284
rect 9852 12282 9858 12299
rect 9829 12279 9858 12282
rect 11967 12278 11970 12304
rect 11996 12298 11999 12304
rect 12106 12299 12135 12302
rect 12106 12298 12112 12299
rect 11996 12284 12112 12298
rect 11996 12278 11999 12284
rect 12106 12282 12112 12284
rect 12129 12282 12135 12299
rect 12574 12298 12588 12347
rect 14313 12346 14316 12372
rect 14342 12346 14345 12372
rect 14322 12332 14336 12346
rect 13540 12318 14336 12332
rect 12795 12298 12798 12304
rect 12574 12284 12798 12298
rect 12106 12279 12135 12282
rect 12795 12278 12798 12284
rect 12824 12298 12827 12304
rect 13540 12298 13554 12318
rect 17211 12312 17214 12338
rect 17240 12332 17243 12338
rect 17266 12332 17280 12376
rect 17312 12366 17326 12420
rect 17671 12380 17674 12406
rect 17700 12400 17703 12406
rect 17764 12401 17793 12404
rect 17764 12400 17770 12401
rect 17700 12386 17770 12400
rect 17700 12380 17703 12386
rect 17764 12384 17770 12386
rect 17787 12400 17793 12401
rect 17818 12400 17832 12454
rect 17864 12420 17970 12434
rect 17864 12406 17878 12420
rect 17787 12386 17832 12400
rect 17787 12384 17793 12386
rect 17764 12381 17793 12384
rect 17855 12380 17858 12406
rect 17884 12380 17887 12406
rect 17901 12380 17904 12406
rect 17930 12380 17933 12406
rect 17956 12400 17970 12420
rect 18315 12414 18318 12440
rect 18344 12414 18347 12440
rect 18416 12438 18430 12454
rect 23974 12452 23980 12469
rect 23997 12468 24003 12469
rect 24249 12468 24252 12474
rect 23997 12454 24252 12468
rect 23997 12452 24003 12454
rect 23974 12449 24003 12452
rect 24249 12448 24252 12454
rect 24278 12448 24281 12474
rect 27147 12448 27150 12474
rect 27176 12448 27179 12474
rect 25583 12438 25586 12440
rect 18408 12435 18437 12438
rect 18408 12418 18414 12435
rect 18431 12418 18437 12435
rect 25565 12435 25586 12438
rect 18408 12415 18437 12418
rect 23890 12420 23996 12434
rect 18454 12401 18483 12404
rect 18454 12400 18460 12401
rect 17956 12386 18460 12400
rect 18454 12384 18460 12386
rect 18477 12384 18483 12401
rect 18454 12381 18483 12384
rect 19143 12380 19146 12406
rect 19172 12380 19175 12406
rect 23890 12404 23904 12420
rect 19236 12401 19265 12404
rect 19236 12400 19242 12401
rect 19198 12386 19242 12400
rect 18591 12366 18594 12372
rect 17312 12352 18594 12366
rect 18591 12346 18594 12352
rect 18620 12366 18623 12372
rect 19198 12366 19212 12386
rect 19236 12384 19242 12386
rect 19259 12384 19265 12401
rect 19236 12381 19265 12384
rect 19282 12401 19311 12404
rect 19282 12384 19288 12401
rect 19305 12384 19311 12401
rect 19282 12381 19311 12384
rect 23882 12401 23911 12404
rect 23882 12384 23888 12401
rect 23905 12384 23911 12401
rect 23882 12381 23911 12384
rect 23928 12401 23957 12404
rect 23928 12384 23934 12401
rect 23951 12384 23957 12401
rect 23982 12400 23996 12420
rect 25565 12418 25571 12435
rect 25565 12415 25586 12418
rect 25583 12414 25586 12415
rect 25612 12414 25615 12440
rect 27331 12414 27334 12440
rect 27360 12414 27363 12440
rect 28113 12414 28116 12440
rect 28142 12434 28145 12440
rect 28274 12435 28303 12438
rect 28274 12434 28280 12435
rect 28142 12420 28280 12434
rect 28142 12414 28145 12420
rect 28274 12418 28280 12420
rect 28297 12418 28303 12435
rect 28274 12415 28303 12418
rect 28325 12435 28354 12438
rect 28325 12418 28331 12435
rect 28348 12434 28354 12435
rect 28389 12434 28392 12440
rect 28348 12420 28392 12434
rect 28348 12418 28354 12420
rect 28325 12415 28354 12418
rect 28389 12414 28392 12420
rect 28418 12414 28421 12440
rect 24433 12400 24436 12406
rect 23982 12386 24436 12400
rect 23928 12381 23957 12384
rect 19290 12366 19304 12381
rect 18620 12352 19212 12366
rect 19244 12352 19304 12366
rect 18620 12346 18623 12352
rect 17240 12318 17280 12332
rect 17240 12312 17243 12318
rect 18315 12312 18318 12338
rect 18344 12332 18347 12338
rect 19244 12332 19258 12352
rect 18344 12318 19258 12332
rect 19282 12333 19311 12336
rect 18344 12312 18347 12318
rect 19282 12316 19288 12333
rect 19305 12332 19311 12333
rect 19373 12332 19376 12338
rect 19305 12318 19376 12332
rect 19305 12316 19311 12318
rect 19282 12313 19311 12316
rect 19373 12312 19376 12318
rect 19402 12312 19405 12338
rect 23936 12332 23950 12381
rect 24433 12380 24436 12386
rect 24462 12380 24465 12406
rect 25354 12401 25383 12404
rect 25354 12384 25360 12401
rect 25377 12400 25383 12401
rect 25399 12400 25402 12406
rect 25377 12386 25402 12400
rect 25377 12384 25383 12386
rect 25354 12381 25383 12384
rect 25399 12380 25402 12386
rect 25428 12380 25431 12406
rect 25515 12401 25544 12404
rect 25515 12384 25521 12401
rect 25538 12400 25544 12401
rect 25629 12400 25632 12406
rect 25538 12386 25632 12400
rect 25538 12384 25544 12386
rect 25515 12381 25544 12384
rect 25629 12380 25632 12386
rect 25658 12380 25661 12406
rect 26389 12401 26418 12404
rect 26389 12384 26395 12401
rect 26412 12400 26418 12401
rect 26642 12401 26671 12404
rect 26642 12400 26648 12401
rect 26412 12386 26648 12400
rect 26412 12384 26418 12386
rect 26389 12381 26418 12384
rect 26642 12384 26648 12386
rect 26665 12384 26671 12401
rect 26642 12381 26671 12384
rect 26687 12380 26690 12406
rect 26716 12400 26719 12406
rect 26734 12401 26763 12404
rect 26734 12400 26740 12401
rect 26716 12386 26740 12400
rect 26716 12380 26719 12386
rect 26734 12384 26740 12386
rect 26757 12384 26763 12401
rect 26734 12381 26763 12384
rect 26779 12380 26782 12406
rect 26808 12380 26811 12406
rect 26826 12401 26855 12404
rect 26826 12384 26832 12401
rect 26849 12400 26855 12401
rect 26871 12400 26874 12406
rect 26849 12386 26874 12400
rect 26849 12384 26855 12386
rect 26826 12381 26855 12384
rect 26871 12380 26874 12386
rect 26900 12380 26903 12406
rect 27148 12401 27177 12404
rect 27148 12400 27154 12401
rect 26926 12386 27154 12400
rect 24065 12346 24068 12372
rect 24094 12346 24097 12372
rect 26926 12336 26940 12386
rect 27148 12384 27154 12386
rect 27171 12384 27177 12401
rect 27148 12381 27177 12384
rect 27193 12380 27196 12406
rect 27222 12380 27225 12406
rect 27286 12401 27315 12404
rect 27286 12384 27292 12401
rect 27309 12384 27315 12401
rect 27286 12381 27315 12384
rect 26918 12333 26947 12336
rect 23936 12318 24732 12332
rect 12824 12284 13554 12298
rect 13601 12299 13630 12302
rect 12824 12278 12827 12284
rect 13601 12282 13607 12299
rect 13624 12298 13630 12299
rect 14221 12298 14224 12304
rect 13624 12284 14224 12298
rect 13624 12282 13630 12284
rect 13601 12279 13630 12282
rect 14221 12278 14224 12284
rect 14250 12278 14253 12304
rect 14911 12278 14914 12304
rect 14940 12298 14943 12304
rect 15349 12299 15378 12302
rect 15349 12298 15355 12299
rect 14940 12284 15355 12298
rect 14940 12278 14943 12284
rect 15349 12282 15355 12284
rect 15372 12282 15378 12299
rect 15349 12279 15378 12282
rect 16291 12278 16294 12304
rect 16320 12278 16323 12304
rect 16981 12278 16984 12304
rect 17010 12298 17013 12304
rect 17074 12299 17103 12302
rect 17074 12298 17080 12299
rect 17010 12284 17080 12298
rect 17010 12278 17013 12284
rect 17074 12282 17080 12284
rect 17097 12282 17103 12299
rect 17074 12279 17103 12282
rect 17533 12278 17536 12304
rect 17562 12298 17565 12304
rect 17810 12299 17839 12302
rect 17810 12298 17816 12299
rect 17562 12284 17816 12298
rect 17562 12278 17565 12284
rect 17810 12282 17816 12284
rect 17833 12282 17839 12299
rect 17810 12279 17839 12282
rect 18454 12299 18483 12302
rect 18454 12282 18460 12299
rect 18477 12298 18483 12299
rect 18499 12298 18502 12304
rect 18477 12284 18502 12298
rect 18477 12282 18483 12284
rect 18454 12279 18483 12282
rect 18499 12278 18502 12284
rect 18528 12278 18531 12304
rect 19419 12278 19422 12304
rect 19448 12298 19451 12304
rect 21489 12298 21492 12304
rect 19448 12284 21492 12298
rect 19448 12278 19451 12284
rect 21489 12278 21492 12284
rect 21518 12278 21521 12304
rect 23927 12278 23930 12304
rect 23956 12278 23959 12304
rect 24718 12298 24732 12318
rect 26918 12316 26924 12333
rect 26941 12316 26947 12333
rect 26918 12313 26947 12316
rect 26825 12298 26828 12304
rect 24718 12284 26828 12298
rect 26825 12278 26828 12284
rect 26854 12278 26857 12304
rect 27294 12298 27308 12381
rect 27377 12380 27380 12406
rect 27406 12380 27409 12406
rect 29149 12401 29178 12404
rect 29149 12384 29155 12401
rect 29172 12400 29178 12401
rect 29677 12400 29680 12406
rect 29172 12386 29680 12400
rect 29172 12384 29178 12386
rect 29149 12381 29178 12384
rect 29677 12380 29680 12386
rect 29706 12380 29709 12406
rect 27837 12346 27840 12372
rect 27866 12366 27869 12372
rect 28113 12366 28116 12372
rect 27866 12352 28116 12366
rect 27866 12346 27869 12352
rect 28113 12346 28116 12352
rect 28142 12346 28145 12372
rect 29585 12298 29588 12304
rect 27294 12284 29588 12298
rect 29585 12278 29588 12284
rect 29614 12278 29617 12304
rect 3036 12216 29992 12264
rect 7413 12176 7416 12202
rect 7442 12176 7445 12202
rect 11209 12197 11238 12200
rect 11209 12180 11215 12197
rect 11232 12196 11238 12197
rect 11553 12196 11556 12202
rect 11232 12182 11556 12196
rect 11232 12180 11238 12182
rect 11209 12177 11238 12180
rect 11553 12176 11556 12182
rect 11582 12176 11585 12202
rect 13991 12176 13994 12202
rect 14020 12196 14023 12202
rect 14222 12197 14251 12200
rect 14222 12196 14228 12197
rect 14020 12182 14228 12196
rect 14020 12176 14023 12182
rect 14222 12180 14228 12182
rect 14245 12180 14251 12197
rect 14222 12177 14251 12180
rect 14681 12176 14684 12202
rect 14710 12196 14713 12202
rect 14866 12197 14895 12200
rect 14866 12196 14872 12197
rect 14710 12182 14872 12196
rect 14710 12176 14713 12182
rect 14866 12180 14872 12182
rect 14889 12180 14895 12197
rect 14866 12177 14895 12180
rect 15693 12176 15696 12202
rect 15722 12196 15725 12202
rect 15786 12197 15815 12200
rect 15786 12196 15792 12197
rect 15722 12182 15792 12196
rect 15722 12176 15725 12182
rect 15786 12180 15792 12182
rect 15809 12180 15815 12197
rect 15786 12177 15815 12180
rect 16797 12176 16800 12202
rect 16826 12196 16829 12202
rect 16982 12197 17011 12200
rect 16982 12196 16988 12197
rect 16826 12182 16988 12196
rect 16826 12176 16829 12182
rect 16982 12180 16988 12182
rect 17005 12180 17011 12197
rect 16982 12177 17011 12180
rect 19143 12176 19146 12202
rect 19172 12196 19175 12202
rect 19926 12197 19955 12200
rect 19926 12196 19932 12197
rect 19172 12182 19932 12196
rect 19172 12176 19175 12182
rect 19926 12180 19932 12182
rect 19949 12180 19955 12197
rect 25399 12196 25402 12202
rect 19926 12177 19955 12180
rect 25224 12182 25402 12196
rect 5389 12142 5392 12168
rect 5418 12162 5421 12168
rect 5574 12163 5603 12166
rect 5574 12162 5580 12163
rect 5418 12148 5580 12162
rect 5418 12142 5421 12148
rect 5574 12146 5580 12148
rect 5597 12146 5603 12163
rect 16107 12162 16110 12168
rect 5574 12143 5603 12146
rect 14460 12148 16110 12162
rect 4515 12108 4518 12134
rect 4544 12128 4547 12134
rect 4700 12129 4729 12132
rect 4700 12128 4706 12129
rect 4544 12114 4706 12128
rect 4544 12108 4547 12114
rect 4700 12112 4706 12114
rect 4723 12128 4729 12129
rect 6839 12129 6868 12132
rect 4723 12114 5826 12128
rect 4723 12112 4729 12114
rect 4700 12109 4729 12112
rect 5812 12098 5826 12114
rect 6839 12112 6845 12129
rect 6862 12128 6868 12129
rect 6862 12114 7620 12128
rect 6862 12112 6868 12114
rect 6839 12109 6868 12112
rect 5804 12095 5833 12098
rect 5804 12078 5810 12095
rect 5827 12094 5833 12095
rect 5849 12094 5852 12100
rect 5827 12080 5852 12094
rect 5827 12078 5833 12080
rect 5804 12075 5833 12078
rect 5849 12074 5852 12080
rect 5878 12074 5881 12100
rect 5941 12074 5944 12100
rect 5970 12098 5973 12100
rect 5970 12095 5988 12098
rect 5982 12078 5988 12095
rect 7321 12094 7324 12100
rect 5970 12075 5988 12078
rect 6134 12080 7324 12094
rect 5970 12074 5973 12075
rect 4837 12040 4840 12066
rect 4866 12040 4869 12066
rect 5527 12060 5530 12066
rect 5451 12046 5530 12060
rect 5527 12040 5530 12046
rect 5556 12060 5559 12066
rect 5665 12060 5668 12066
rect 5556 12046 5668 12060
rect 5556 12040 5559 12046
rect 5665 12040 5668 12046
rect 5694 12040 5697 12066
rect 6015 12061 6044 12064
rect 6015 12044 6021 12061
rect 6038 12060 6044 12061
rect 6134 12060 6148 12080
rect 7321 12074 7324 12080
rect 7350 12074 7353 12100
rect 7413 12074 7416 12100
rect 7442 12074 7445 12100
rect 7459 12074 7462 12100
rect 7488 12074 7491 12100
rect 7551 12074 7554 12100
rect 7580 12074 7583 12100
rect 7606 12098 7620 12114
rect 8471 12108 8474 12134
rect 8500 12128 8503 12134
rect 8522 12129 8551 12132
rect 8522 12128 8528 12129
rect 8500 12114 8528 12128
rect 8500 12108 8503 12114
rect 8522 12112 8528 12114
rect 8545 12112 8551 12129
rect 8522 12109 8551 12112
rect 10035 12108 10038 12134
rect 10064 12128 10067 12134
rect 10174 12129 10203 12132
rect 10174 12128 10180 12129
rect 10064 12114 10180 12128
rect 10064 12108 10067 12114
rect 10174 12112 10180 12114
rect 10197 12112 10203 12129
rect 10174 12109 10203 12112
rect 11967 12108 11970 12134
rect 11996 12108 11999 12134
rect 13853 12108 13856 12134
rect 13882 12128 13885 12134
rect 13882 12114 14336 12128
rect 13882 12108 13885 12114
rect 7598 12095 7627 12098
rect 7598 12078 7604 12095
rect 7621 12078 7627 12095
rect 7598 12075 7627 12078
rect 7644 12095 7673 12098
rect 7644 12078 7650 12095
rect 7667 12094 7673 12095
rect 9115 12094 9118 12100
rect 7667 12080 9118 12094
rect 7667 12078 7673 12080
rect 7644 12075 7673 12078
rect 9115 12074 9118 12080
rect 9144 12074 9147 12100
rect 10219 12074 10222 12100
rect 10248 12094 10251 12100
rect 10335 12095 10364 12098
rect 10335 12094 10341 12095
rect 10248 12080 10341 12094
rect 10248 12074 10251 12080
rect 10335 12078 10341 12080
rect 10358 12094 10364 12095
rect 10449 12094 10452 12100
rect 10358 12080 10452 12094
rect 10358 12078 10364 12080
rect 10335 12075 10364 12078
rect 10449 12074 10452 12080
rect 10478 12074 10481 12100
rect 12013 12074 12016 12100
rect 12042 12098 12045 12100
rect 12042 12094 12046 12098
rect 12042 12080 12064 12094
rect 12042 12075 12046 12080
rect 12042 12074 12045 12075
rect 12795 12074 12798 12100
rect 12824 12094 12827 12100
rect 12934 12095 12963 12098
rect 12934 12094 12940 12095
rect 12824 12080 12940 12094
rect 12824 12074 12827 12080
rect 12934 12078 12940 12080
rect 12957 12078 12963 12095
rect 12934 12075 12963 12078
rect 14221 12074 14224 12100
rect 14250 12074 14253 12100
rect 14322 12098 14336 12114
rect 14314 12095 14343 12098
rect 14314 12078 14320 12095
rect 14337 12078 14343 12095
rect 14314 12075 14343 12078
rect 14405 12074 14408 12100
rect 14434 12098 14437 12100
rect 14434 12094 14438 12098
rect 14460 12094 14474 12148
rect 16107 12142 16110 12148
rect 16136 12142 16139 12168
rect 19281 12162 19284 12168
rect 17404 12148 19284 12162
rect 16223 12129 16252 12132
rect 16223 12128 16229 12129
rect 15932 12114 16229 12128
rect 15932 12100 15946 12114
rect 16223 12112 16229 12114
rect 16246 12112 16252 12129
rect 16223 12109 16252 12112
rect 14434 12080 14474 12094
rect 14434 12075 14438 12080
rect 14434 12074 14437 12075
rect 14819 12074 14822 12100
rect 14848 12074 14851 12100
rect 14911 12074 14914 12100
rect 14940 12074 14943 12100
rect 15923 12074 15926 12100
rect 15952 12074 15955 12100
rect 16107 12074 16110 12100
rect 16136 12094 16139 12100
rect 16172 12095 16201 12098
rect 16172 12094 16178 12095
rect 16136 12080 16178 12094
rect 16136 12074 16139 12080
rect 16172 12078 16178 12080
rect 16195 12078 16201 12095
rect 16172 12075 16201 12078
rect 16981 12074 16984 12100
rect 17010 12074 17013 12100
rect 17074 12095 17103 12098
rect 17074 12078 17080 12095
rect 17097 12078 17103 12095
rect 17074 12075 17103 12078
rect 6038 12046 6148 12060
rect 6038 12044 6044 12046
rect 6015 12041 6044 12044
rect 8563 12040 8566 12066
rect 8592 12060 8595 12066
rect 8678 12061 8707 12064
rect 8678 12060 8684 12061
rect 8592 12046 8684 12060
rect 8592 12040 8595 12046
rect 8678 12044 8684 12046
rect 8701 12044 8707 12061
rect 8678 12041 8707 12044
rect 8729 12061 8758 12064
rect 8729 12044 8735 12061
rect 8752 12060 8758 12061
rect 8793 12060 8796 12066
rect 8752 12046 8796 12060
rect 8752 12044 8758 12046
rect 8729 12041 8758 12044
rect 8793 12040 8796 12046
rect 8822 12040 8825 12066
rect 10403 12064 10406 12066
rect 10385 12061 10406 12064
rect 10385 12044 10391 12061
rect 10385 12041 10406 12044
rect 10403 12040 10406 12041
rect 10432 12040 10435 12066
rect 11829 12040 11832 12066
rect 11858 12040 11861 12066
rect 11921 12040 11924 12066
rect 11950 12040 11953 12066
rect 11967 12040 11970 12066
rect 11996 12040 11999 12066
rect 12887 12040 12890 12066
rect 12916 12060 12919 12066
rect 13163 12064 13166 12066
rect 13094 12061 13123 12064
rect 13094 12060 13100 12061
rect 12916 12046 13100 12060
rect 12916 12040 12919 12046
rect 13094 12044 13100 12046
rect 13117 12044 13123 12061
rect 13094 12041 13123 12044
rect 13145 12061 13166 12064
rect 13145 12044 13151 12061
rect 13145 12041 13166 12044
rect 13163 12040 13166 12041
rect 13192 12040 13195 12066
rect 14360 12061 14389 12064
rect 14360 12044 14366 12061
rect 14383 12044 14389 12061
rect 14360 12041 14389 12044
rect 9529 12006 9532 12032
rect 9558 12030 9561 12032
rect 9558 12027 9582 12030
rect 9558 12010 9559 12027
rect 9576 12010 9582 12027
rect 9558 12007 9582 12010
rect 13969 12027 13998 12030
rect 13969 12010 13975 12027
rect 13992 12026 13998 12027
rect 14368 12026 14382 12041
rect 15785 12040 15788 12066
rect 15814 12040 15817 12066
rect 15878 12061 15907 12064
rect 15878 12044 15884 12061
rect 15901 12060 15907 12061
rect 16291 12060 16294 12066
rect 15901 12046 16294 12060
rect 15901 12044 15907 12046
rect 15878 12041 15907 12044
rect 16291 12040 16294 12046
rect 16320 12040 16323 12066
rect 16567 12040 16570 12066
rect 16596 12060 16599 12066
rect 17082 12060 17096 12075
rect 17257 12074 17260 12100
rect 17286 12094 17289 12100
rect 17404 12098 17418 12148
rect 19281 12142 19284 12148
rect 19310 12142 19313 12168
rect 19511 12142 19514 12168
rect 19540 12142 19543 12168
rect 21996 12163 22025 12166
rect 21996 12162 22002 12163
rect 19842 12148 22002 12162
rect 18499 12108 18502 12134
rect 18528 12108 18531 12134
rect 18637 12108 18640 12134
rect 18666 12128 18669 12134
rect 18730 12129 18759 12132
rect 18730 12128 18736 12129
rect 18666 12114 18736 12128
rect 18666 12108 18669 12114
rect 18730 12112 18736 12114
rect 18753 12112 18759 12129
rect 18730 12109 18759 12112
rect 17396 12095 17425 12098
rect 17396 12094 17402 12095
rect 17286 12080 17402 12094
rect 17286 12074 17289 12080
rect 17396 12078 17402 12080
rect 17419 12078 17425 12095
rect 17396 12075 17425 12078
rect 17533 12074 17536 12100
rect 17562 12074 17565 12100
rect 17901 12074 17904 12100
rect 17930 12094 17933 12100
rect 18546 12095 18575 12098
rect 18546 12094 18552 12095
rect 17930 12080 18552 12094
rect 17930 12074 17933 12080
rect 18546 12078 18552 12080
rect 18569 12078 18575 12095
rect 19290 12094 19304 12142
rect 19842 12132 19856 12148
rect 21996 12146 22002 12148
rect 22019 12146 22025 12163
rect 21996 12143 22025 12146
rect 19834 12129 19863 12132
rect 19834 12112 19840 12129
rect 19857 12112 19863 12129
rect 19834 12109 19863 12112
rect 19972 12129 20001 12132
rect 19972 12112 19978 12129
rect 19995 12112 20001 12129
rect 22593 12128 22596 12134
rect 19972 12109 20001 12112
rect 21958 12114 22596 12128
rect 19466 12095 19495 12098
rect 19466 12094 19472 12095
rect 19290 12080 19472 12094
rect 18546 12075 18575 12078
rect 19466 12078 19472 12080
rect 19489 12078 19495 12095
rect 19466 12075 19495 12078
rect 16596 12046 17096 12060
rect 18554 12060 18568 12075
rect 19879 12074 19882 12100
rect 19908 12074 19911 12100
rect 19373 12060 19376 12066
rect 18554 12046 19376 12060
rect 16596 12040 16599 12046
rect 19373 12040 19376 12046
rect 19402 12060 19405 12066
rect 19604 12061 19633 12064
rect 19604 12060 19610 12061
rect 19402 12046 19610 12060
rect 19402 12040 19405 12046
rect 19604 12044 19610 12046
rect 19627 12044 19633 12061
rect 19980 12060 19994 12109
rect 21958 12098 21972 12114
rect 22593 12108 22596 12114
rect 22622 12108 22625 12134
rect 25224 12132 25238 12182
rect 25399 12176 25402 12182
rect 25428 12176 25431 12202
rect 26251 12197 26280 12200
rect 26251 12180 26257 12197
rect 26274 12196 26280 12197
rect 26779 12196 26782 12202
rect 26274 12182 26782 12196
rect 26274 12180 26280 12182
rect 26251 12177 26280 12180
rect 26779 12176 26782 12182
rect 26808 12176 26811 12202
rect 25216 12129 25245 12132
rect 25216 12112 25222 12129
rect 25239 12112 25245 12129
rect 25216 12109 25245 12112
rect 21950 12095 21979 12098
rect 21950 12078 21956 12095
rect 21973 12078 21979 12095
rect 21950 12075 21979 12078
rect 22087 12074 22090 12100
rect 22116 12074 22119 12100
rect 25377 12095 25406 12098
rect 25377 12078 25383 12095
rect 25400 12094 25406 12095
rect 25629 12094 25632 12100
rect 25400 12080 25632 12094
rect 25400 12078 25406 12080
rect 25377 12075 25406 12078
rect 25629 12074 25632 12080
rect 25658 12074 25661 12100
rect 19604 12041 19633 12044
rect 19658 12046 19994 12060
rect 13992 12012 14382 12026
rect 13992 12010 13998 12012
rect 13969 12007 13998 12010
rect 9558 12006 9561 12007
rect 16659 12006 16662 12032
rect 16688 12026 16691 12032
rect 17165 12026 17168 12032
rect 16688 12012 17168 12026
rect 16688 12006 16691 12012
rect 17165 12006 17168 12012
rect 17194 12026 17197 12032
rect 17442 12027 17471 12030
rect 17442 12026 17448 12027
rect 17194 12012 17448 12026
rect 17194 12006 17197 12012
rect 17442 12010 17448 12012
rect 17465 12010 17471 12027
rect 17442 12007 17471 12010
rect 19465 12006 19468 12032
rect 19494 12026 19497 12032
rect 19658 12026 19672 12046
rect 21581 12040 21584 12066
rect 21610 12060 21613 12066
rect 22042 12061 22071 12064
rect 22042 12060 22048 12061
rect 21610 12046 22048 12060
rect 21610 12040 21613 12046
rect 22042 12044 22048 12046
rect 22065 12044 22071 12061
rect 22042 12041 22071 12044
rect 25427 12061 25456 12064
rect 25427 12044 25433 12061
rect 25450 12060 25456 12061
rect 25491 12060 25494 12066
rect 25450 12046 25494 12060
rect 25450 12044 25456 12046
rect 25427 12041 25456 12044
rect 25491 12040 25494 12046
rect 25520 12040 25523 12066
rect 19494 12012 19672 12026
rect 19494 12006 19497 12012
rect 3036 11944 29992 11992
rect 4837 11904 4840 11930
rect 4866 11924 4869 11930
rect 5206 11925 5235 11928
rect 5206 11924 5212 11925
rect 4866 11910 5212 11924
rect 4866 11904 4869 11910
rect 5206 11908 5212 11910
rect 5229 11908 5235 11925
rect 5206 11905 5235 11908
rect 5389 11904 5392 11930
rect 5418 11904 5421 11930
rect 5435 11904 5438 11930
rect 5464 11904 5467 11930
rect 9208 11925 9237 11928
rect 9208 11908 9214 11925
rect 9231 11908 9237 11925
rect 9208 11905 9237 11908
rect 10979 11925 11008 11928
rect 10979 11908 10985 11925
rect 11002 11924 11008 11925
rect 11691 11924 11694 11930
rect 11002 11910 11694 11924
rect 11002 11908 11008 11910
rect 10979 11905 11008 11908
rect 7321 11870 7324 11896
rect 7350 11890 7353 11896
rect 7483 11891 7512 11894
rect 7483 11890 7489 11891
rect 7350 11876 7489 11890
rect 7350 11870 7353 11876
rect 7483 11874 7489 11876
rect 7506 11874 7512 11891
rect 7483 11871 7512 11874
rect 8311 11891 8340 11894
rect 8311 11874 8317 11891
rect 8334 11890 8340 11891
rect 9070 11891 9099 11894
rect 9070 11890 9076 11891
rect 8334 11876 9076 11890
rect 8334 11874 8340 11876
rect 8311 11871 8340 11874
rect 9070 11874 9076 11876
rect 9093 11874 9099 11891
rect 9070 11871 9099 11874
rect 5895 11836 5898 11862
rect 5924 11856 5927 11862
rect 6080 11857 6109 11860
rect 6080 11856 6086 11857
rect 5924 11842 6086 11856
rect 5924 11836 5927 11842
rect 6080 11840 6086 11842
rect 6103 11840 6109 11857
rect 6080 11837 6109 11840
rect 7091 11836 7094 11862
rect 7120 11856 7123 11862
rect 7437 11857 7466 11860
rect 7437 11856 7443 11857
rect 7120 11842 7443 11856
rect 7120 11836 7123 11842
rect 7437 11840 7443 11842
rect 7460 11856 7466 11857
rect 8609 11856 8612 11862
rect 7460 11842 8612 11856
rect 7460 11840 7466 11842
rect 7437 11837 7466 11840
rect 8609 11836 8612 11842
rect 8638 11836 8641 11862
rect 8931 11836 8934 11862
rect 8960 11836 8963 11862
rect 8977 11836 8980 11862
rect 9006 11856 9009 11862
rect 9024 11857 9053 11860
rect 9024 11856 9030 11857
rect 9006 11842 9030 11856
rect 9006 11836 9009 11842
rect 9024 11840 9030 11842
rect 9047 11840 9053 11857
rect 9024 11837 9053 11840
rect 9115 11836 9118 11862
rect 9144 11836 9147 11862
rect 9216 11856 9230 11905
rect 11691 11904 11694 11910
rect 11720 11904 11723 11930
rect 15785 11904 15788 11930
rect 15814 11924 15817 11930
rect 16108 11925 16137 11928
rect 16108 11924 16114 11925
rect 15814 11910 16114 11924
rect 15814 11904 15817 11910
rect 16108 11908 16114 11910
rect 16131 11908 16137 11925
rect 16108 11905 16137 11908
rect 19373 11904 19376 11930
rect 19402 11904 19405 11930
rect 26941 11925 26970 11928
rect 26941 11908 26947 11925
rect 26964 11924 26970 11925
rect 27193 11924 27196 11930
rect 26964 11910 27196 11924
rect 26964 11908 26970 11910
rect 26941 11905 26970 11908
rect 27193 11904 27196 11910
rect 27222 11904 27225 11930
rect 9622 11891 9651 11894
rect 9622 11874 9628 11891
rect 9645 11890 9651 11891
rect 9713 11890 9716 11896
rect 9645 11876 9716 11890
rect 9645 11874 9651 11876
rect 9622 11871 9651 11874
rect 9713 11870 9716 11876
rect 9742 11870 9745 11896
rect 9989 11870 9992 11896
rect 10018 11890 10021 11896
rect 13025 11894 13028 11896
rect 10151 11891 10180 11894
rect 10151 11890 10157 11891
rect 10018 11876 10157 11890
rect 10018 11870 10021 11876
rect 10151 11874 10157 11876
rect 10174 11890 10180 11891
rect 13007 11891 13028 11894
rect 10174 11876 10288 11890
rect 10174 11874 10180 11876
rect 10151 11871 10180 11874
rect 9438 11857 9467 11860
rect 9438 11856 9444 11857
rect 9216 11842 9444 11856
rect 9438 11840 9444 11842
rect 9461 11840 9467 11857
rect 9438 11837 9467 11840
rect 9484 11857 9513 11860
rect 9484 11840 9490 11857
rect 9507 11856 9513 11857
rect 9529 11856 9532 11862
rect 9507 11842 9532 11856
rect 9507 11840 9513 11842
rect 9484 11837 9513 11840
rect 9529 11836 9532 11842
rect 9558 11836 9561 11862
rect 9575 11836 9578 11862
rect 9604 11836 9607 11862
rect 9667 11836 9670 11862
rect 9696 11836 9699 11862
rect 10105 11857 10134 11860
rect 10105 11840 10111 11857
rect 10128 11856 10134 11857
rect 10219 11856 10222 11862
rect 10128 11842 10222 11856
rect 10128 11840 10134 11842
rect 10105 11837 10134 11840
rect 10219 11836 10222 11842
rect 10248 11836 10251 11862
rect 10274 11856 10288 11876
rect 13007 11874 13013 11891
rect 13007 11871 13028 11874
rect 13025 11870 13028 11871
rect 13054 11870 13057 11896
rect 13831 11891 13860 11894
rect 13831 11874 13837 11891
rect 13854 11890 13860 11891
rect 14452 11891 14481 11894
rect 14452 11890 14458 11891
rect 13854 11876 14458 11890
rect 13854 11874 13860 11876
rect 13831 11871 13860 11874
rect 14452 11874 14458 11876
rect 14475 11874 14481 11891
rect 16383 11890 16386 11896
rect 14452 11871 14481 11874
rect 16116 11876 16386 11890
rect 11876 11857 11905 11860
rect 10274 11842 10840 11856
rect 5343 11802 5346 11828
rect 5372 11822 5375 11828
rect 5481 11822 5484 11828
rect 5372 11808 5484 11822
rect 5372 11802 5375 11808
rect 5481 11802 5484 11808
rect 5510 11802 5513 11828
rect 6861 11802 6864 11828
rect 6890 11802 6893 11828
rect 7046 11823 7075 11826
rect 7046 11806 7052 11823
rect 7069 11822 7075 11823
rect 7276 11823 7305 11826
rect 7276 11822 7282 11823
rect 7069 11808 7282 11822
rect 7069 11806 7075 11808
rect 7046 11803 7075 11806
rect 7276 11806 7282 11808
rect 7299 11806 7305 11823
rect 7276 11803 7305 11806
rect 9714 11823 9743 11826
rect 9714 11806 9720 11823
rect 9737 11822 9743 11823
rect 9897 11822 9900 11828
rect 9737 11808 9900 11822
rect 9737 11806 9743 11808
rect 9714 11803 9743 11806
rect 9897 11802 9900 11808
rect 9926 11802 9929 11828
rect 9944 11823 9973 11826
rect 9944 11806 9950 11823
rect 9967 11806 9973 11823
rect 9944 11803 9973 11806
rect 9952 11754 9966 11803
rect 10826 11788 10840 11842
rect 11876 11840 11882 11857
rect 11899 11856 11905 11857
rect 12795 11856 12798 11862
rect 11899 11842 12798 11856
rect 11899 11840 11905 11842
rect 11876 11837 11905 11840
rect 10863 11802 10866 11828
rect 10892 11822 10895 11828
rect 11884 11822 11898 11837
rect 12795 11836 12798 11842
rect 12824 11836 12827 11862
rect 12933 11836 12936 11862
rect 12962 11860 12965 11862
rect 12962 11857 12980 11860
rect 12974 11840 12980 11857
rect 12962 11837 12980 11840
rect 12962 11836 12965 11837
rect 14313 11836 14316 11862
rect 14342 11836 14345 11862
rect 14359 11836 14362 11862
rect 14388 11856 14391 11862
rect 14406 11857 14435 11860
rect 14406 11856 14412 11857
rect 14388 11842 14412 11856
rect 14388 11836 14391 11842
rect 14406 11840 14412 11842
rect 14429 11840 14435 11857
rect 14406 11837 14435 11840
rect 14497 11836 14500 11862
rect 14526 11860 14529 11862
rect 14526 11856 14530 11860
rect 15969 11856 15972 11862
rect 14526 11842 15972 11856
rect 14526 11837 14530 11842
rect 14526 11836 14529 11837
rect 15969 11836 15972 11842
rect 15998 11836 16001 11862
rect 16116 11860 16130 11876
rect 16383 11870 16386 11876
rect 16412 11870 16415 11896
rect 20413 11891 20442 11894
rect 18692 11876 19327 11890
rect 16108 11857 16137 11860
rect 16108 11840 16114 11857
rect 16131 11840 16137 11857
rect 16108 11837 16137 11840
rect 16245 11836 16248 11862
rect 16274 11836 16277 11862
rect 16292 11857 16321 11860
rect 16292 11840 16298 11857
rect 16315 11856 16321 11857
rect 16337 11856 16340 11862
rect 16315 11842 16340 11856
rect 16315 11840 16321 11842
rect 16292 11837 16321 11840
rect 16337 11836 16340 11842
rect 16366 11856 16369 11862
rect 16521 11856 16524 11862
rect 16366 11842 16524 11856
rect 16366 11836 16369 11842
rect 16521 11836 16524 11842
rect 16550 11836 16553 11862
rect 18692 11860 18706 11876
rect 18684 11857 18713 11860
rect 18684 11840 18690 11857
rect 18707 11840 18713 11857
rect 18684 11837 18713 11840
rect 18729 11836 18732 11862
rect 18758 11856 18761 11862
rect 18812 11857 18841 11860
rect 18812 11856 18818 11857
rect 18758 11842 18818 11856
rect 18758 11836 18761 11842
rect 18812 11840 18818 11842
rect 18835 11840 18841 11857
rect 18812 11837 18841 11840
rect 10892 11808 11898 11822
rect 10892 11802 10895 11808
rect 12381 11802 12384 11828
rect 12410 11802 12413 11828
rect 19313 11822 19327 11876
rect 20413 11874 20419 11891
rect 20436 11890 20442 11891
rect 20436 11876 20546 11890
rect 20436 11874 20442 11876
rect 20413 11871 20442 11874
rect 20109 11836 20112 11862
rect 20138 11856 20141 11862
rect 20357 11857 20386 11860
rect 20357 11856 20363 11857
rect 20138 11842 20363 11856
rect 20138 11836 20141 11842
rect 20357 11840 20363 11842
rect 20380 11856 20386 11857
rect 20477 11856 20480 11862
rect 20380 11842 20480 11856
rect 20380 11840 20386 11842
rect 20357 11837 20386 11840
rect 20477 11836 20480 11842
rect 20506 11836 20509 11862
rect 20532 11856 20546 11876
rect 21443 11870 21446 11896
rect 21472 11890 21475 11896
rect 21472 11876 21650 11890
rect 21472 11870 21475 11876
rect 21636 11862 21650 11876
rect 25629 11870 25632 11896
rect 25658 11890 25661 11896
rect 26066 11891 26095 11894
rect 26066 11890 26072 11891
rect 25658 11876 26072 11890
rect 25658 11870 25661 11876
rect 26066 11874 26072 11876
rect 26089 11874 26095 11891
rect 26066 11871 26095 11874
rect 26117 11891 26146 11894
rect 26117 11874 26123 11891
rect 26140 11890 26146 11891
rect 26181 11890 26184 11896
rect 26140 11876 26184 11890
rect 26140 11874 26146 11876
rect 26117 11871 26146 11874
rect 26181 11870 26184 11876
rect 26210 11870 26213 11896
rect 20753 11856 20756 11862
rect 20532 11842 20756 11856
rect 20753 11836 20756 11842
rect 20782 11856 20785 11862
rect 20845 11856 20848 11862
rect 20782 11842 20848 11856
rect 20782 11836 20785 11842
rect 20845 11836 20848 11842
rect 20874 11836 20877 11862
rect 21237 11857 21266 11860
rect 21237 11840 21243 11857
rect 21260 11856 21266 11857
rect 21536 11857 21565 11860
rect 21536 11856 21542 11857
rect 21260 11842 21542 11856
rect 21260 11840 21266 11842
rect 21237 11837 21266 11840
rect 21536 11840 21542 11842
rect 21559 11840 21565 11857
rect 21536 11837 21565 11840
rect 21627 11836 21630 11862
rect 21656 11836 21659 11862
rect 21673 11836 21676 11862
rect 21702 11836 21705 11862
rect 21719 11836 21722 11862
rect 21748 11860 21751 11862
rect 21748 11856 21752 11860
rect 21748 11842 21770 11856
rect 21748 11837 21752 11842
rect 21748 11836 21751 11837
rect 25399 11836 25402 11862
rect 25428 11856 25431 11862
rect 25906 11857 25935 11860
rect 25906 11856 25912 11857
rect 25428 11842 25912 11856
rect 25428 11836 25431 11842
rect 25906 11840 25912 11842
rect 25929 11840 25935 11857
rect 25906 11837 25935 11840
rect 20155 11822 20158 11828
rect 19313 11808 20158 11822
rect 20155 11802 20158 11808
rect 20184 11822 20187 11828
rect 20202 11823 20231 11826
rect 20202 11822 20208 11823
rect 20184 11808 20208 11822
rect 20184 11802 20187 11808
rect 20202 11806 20208 11808
rect 20225 11806 20231 11823
rect 20202 11803 20231 11806
rect 21581 11802 21584 11828
rect 21610 11802 21613 11828
rect 10826 11774 11047 11788
rect 10863 11754 10866 11760
rect 9952 11740 10866 11754
rect 10863 11734 10866 11740
rect 10892 11734 10895 11760
rect 11033 11754 11047 11774
rect 14037 11768 14040 11794
rect 14066 11788 14069 11794
rect 14314 11789 14343 11792
rect 14314 11788 14320 11789
rect 14066 11774 14320 11788
rect 14066 11768 14069 11774
rect 14314 11772 14320 11774
rect 14337 11772 14343 11789
rect 14314 11769 14343 11772
rect 13163 11754 13166 11760
rect 11033 11740 13166 11754
rect 13163 11734 13166 11740
rect 13192 11734 13195 11760
rect 19925 11734 19928 11760
rect 19954 11754 19957 11760
rect 21719 11754 21722 11760
rect 19954 11740 21722 11754
rect 19954 11734 19957 11740
rect 21719 11734 21722 11740
rect 21748 11734 21751 11760
rect 3036 11672 29992 11720
rect 7413 11632 7416 11658
rect 7442 11652 7445 11658
rect 7690 11653 7719 11656
rect 7690 11652 7696 11653
rect 7442 11638 7696 11652
rect 7442 11632 7445 11638
rect 7690 11636 7696 11638
rect 7713 11636 7719 11653
rect 9575 11652 9578 11658
rect 7690 11633 7719 11636
rect 8664 11638 9578 11652
rect 8664 11618 8678 11638
rect 9575 11632 9578 11638
rect 9604 11632 9607 11658
rect 9713 11656 9716 11658
rect 9691 11653 9716 11656
rect 9691 11636 9697 11653
rect 9714 11636 9716 11653
rect 9691 11633 9716 11636
rect 9713 11632 9716 11633
rect 9742 11632 9745 11658
rect 11645 11632 11648 11658
rect 11674 11652 11677 11658
rect 11674 11638 11806 11652
rect 11674 11632 11677 11638
rect 7514 11604 8678 11618
rect 11792 11618 11806 11638
rect 11967 11632 11970 11658
rect 11996 11656 11999 11658
rect 11996 11653 12020 11656
rect 11996 11636 11997 11653
rect 12014 11636 12020 11653
rect 13071 11652 13074 11658
rect 11996 11633 12020 11636
rect 12068 11638 13074 11652
rect 11996 11632 11999 11633
rect 12068 11618 12082 11638
rect 13071 11632 13074 11638
rect 13100 11632 13103 11658
rect 13969 11653 13998 11656
rect 13969 11636 13975 11653
rect 13992 11652 13998 11653
rect 14313 11652 14316 11658
rect 13992 11638 14316 11652
rect 13992 11636 13998 11638
rect 13969 11633 13998 11636
rect 14313 11632 14316 11638
rect 14342 11632 14345 11658
rect 18684 11653 18713 11656
rect 18684 11636 18690 11653
rect 18707 11652 18713 11653
rect 18729 11652 18732 11658
rect 18707 11638 18732 11652
rect 18707 11636 18713 11638
rect 18684 11633 18713 11636
rect 18729 11632 18732 11638
rect 18758 11632 18761 11658
rect 11792 11604 12082 11618
rect 5895 11530 5898 11556
rect 5924 11530 5927 11556
rect 5941 11530 5944 11556
rect 5970 11550 5973 11556
rect 6057 11551 6086 11554
rect 6057 11550 6063 11551
rect 5970 11536 6063 11550
rect 5970 11530 5973 11536
rect 6057 11534 6063 11536
rect 6080 11550 6086 11551
rect 6171 11550 6174 11556
rect 6080 11536 6174 11550
rect 6080 11534 6086 11536
rect 6057 11531 6086 11534
rect 6171 11530 6174 11536
rect 6200 11530 6203 11556
rect 7514 11554 7528 11604
rect 8471 11564 8474 11590
rect 8500 11584 8503 11590
rect 8656 11585 8685 11588
rect 8656 11584 8662 11585
rect 8500 11570 8662 11584
rect 8500 11564 8503 11570
rect 8656 11568 8662 11570
rect 8679 11568 8685 11585
rect 8656 11565 8685 11568
rect 10173 11564 10176 11590
rect 10202 11584 10205 11590
rect 10202 11570 10334 11584
rect 10202 11564 10205 11570
rect 6931 11551 6960 11554
rect 6931 11534 6937 11551
rect 6954 11550 6960 11551
rect 7414 11551 7443 11554
rect 7414 11550 7420 11551
rect 6954 11536 7420 11550
rect 6954 11534 6960 11536
rect 6931 11531 6960 11534
rect 7414 11534 7420 11536
rect 7437 11534 7443 11551
rect 7414 11531 7443 11534
rect 7506 11551 7535 11554
rect 7506 11534 7512 11551
rect 7529 11534 7535 11551
rect 7506 11531 7535 11534
rect 7597 11530 7600 11556
rect 7626 11530 7629 11556
rect 8701 11530 8704 11556
rect 8730 11550 8733 11556
rect 8855 11551 8884 11554
rect 8855 11550 8861 11551
rect 8730 11536 8861 11550
rect 8730 11530 8733 11536
rect 8855 11534 8861 11536
rect 8878 11550 8884 11551
rect 8878 11536 9690 11550
rect 8878 11534 8884 11536
rect 8855 11531 8884 11534
rect 6125 11520 6128 11522
rect 6107 11517 6128 11520
rect 6107 11500 6113 11517
rect 6107 11497 6128 11500
rect 6125 11496 6128 11497
rect 6154 11496 6157 11522
rect 7551 11496 7554 11522
rect 7580 11496 7583 11522
rect 8609 11496 8612 11522
rect 8638 11516 8641 11522
rect 8816 11517 8845 11520
rect 8816 11516 8822 11517
rect 8638 11502 8822 11516
rect 8638 11496 8641 11502
rect 8816 11500 8822 11502
rect 8839 11500 8845 11517
rect 8816 11497 8845 11500
rect 9676 11482 9690 11536
rect 9897 11530 9900 11556
rect 9926 11550 9929 11556
rect 10320 11554 10334 11570
rect 10449 11564 10452 11590
rect 10478 11584 10481 11590
rect 10478 11570 11024 11584
rect 10478 11564 10481 11570
rect 10266 11551 10295 11554
rect 10266 11550 10272 11551
rect 9926 11536 10272 11550
rect 9926 11530 9929 11536
rect 10266 11534 10272 11536
rect 10289 11534 10295 11551
rect 10266 11531 10295 11534
rect 10312 11551 10341 11554
rect 10312 11534 10318 11551
rect 10335 11534 10341 11551
rect 10312 11531 10341 11534
rect 10863 11530 10866 11556
rect 10892 11550 10895 11556
rect 10956 11551 10985 11554
rect 10956 11550 10962 11551
rect 10892 11536 10962 11550
rect 10892 11530 10895 11536
rect 10956 11534 10962 11536
rect 10979 11534 10985 11551
rect 11010 11550 11024 11570
rect 12795 11564 12798 11590
rect 12824 11584 12827 11590
rect 12934 11585 12963 11588
rect 12934 11584 12940 11585
rect 12824 11570 12940 11584
rect 12824 11564 12827 11570
rect 12934 11568 12940 11570
rect 12957 11568 12963 11585
rect 12934 11565 12963 11568
rect 16476 11585 16505 11588
rect 16476 11568 16482 11585
rect 16499 11584 16505 11585
rect 16659 11584 16662 11590
rect 16499 11570 16662 11584
rect 16499 11568 16505 11570
rect 16476 11565 16505 11568
rect 16659 11564 16662 11570
rect 16688 11564 16691 11590
rect 17441 11564 17444 11590
rect 17470 11584 17473 11590
rect 21167 11584 21170 11590
rect 17470 11570 21170 11584
rect 17470 11564 17473 11570
rect 21167 11564 21170 11570
rect 21196 11564 21199 11590
rect 11093 11550 11096 11556
rect 11122 11554 11125 11556
rect 11122 11551 11140 11554
rect 11010 11536 11096 11550
rect 10956 11531 10985 11534
rect 11093 11530 11096 11536
rect 11134 11534 11140 11551
rect 12979 11550 12982 11556
rect 11122 11531 11140 11534
rect 11286 11536 12982 11550
rect 11122 11530 11125 11531
rect 9943 11496 9946 11522
rect 9972 11516 9975 11522
rect 10174 11517 10203 11520
rect 10174 11516 10180 11517
rect 9972 11502 10180 11516
rect 9972 11496 9975 11502
rect 10174 11500 10180 11502
rect 10197 11500 10203 11517
rect 11167 11517 11196 11520
rect 11167 11516 11173 11517
rect 10174 11497 10203 11500
rect 10228 11502 11173 11516
rect 10228 11482 10242 11502
rect 11167 11500 11173 11502
rect 11190 11516 11196 11517
rect 11286 11516 11300 11536
rect 12979 11530 12982 11536
rect 13008 11530 13011 11556
rect 16337 11530 16340 11556
rect 16366 11530 16369 11556
rect 16383 11530 16386 11556
rect 16412 11530 16415 11556
rect 18637 11530 18640 11556
rect 18666 11530 18669 11556
rect 18729 11530 18732 11556
rect 18758 11530 18761 11556
rect 19465 11530 19468 11556
rect 19494 11530 19497 11556
rect 19558 11551 19587 11554
rect 19558 11534 19564 11551
rect 19581 11550 19587 11551
rect 19833 11550 19836 11556
rect 19581 11536 19836 11550
rect 19581 11534 19587 11536
rect 19558 11531 19587 11534
rect 19833 11530 19836 11536
rect 19862 11550 19865 11556
rect 19925 11550 19928 11556
rect 19862 11536 19928 11550
rect 19862 11530 19865 11536
rect 19925 11530 19928 11536
rect 19954 11530 19957 11556
rect 11190 11502 11300 11516
rect 11190 11500 11196 11502
rect 11167 11497 11196 11500
rect 12933 11496 12936 11522
rect 12962 11516 12965 11522
rect 13163 11520 13166 11522
rect 13094 11517 13123 11520
rect 13094 11516 13100 11517
rect 12962 11502 13100 11516
rect 12962 11496 12965 11502
rect 13094 11500 13100 11502
rect 13117 11500 13123 11517
rect 13094 11497 13123 11500
rect 13145 11517 13166 11520
rect 13145 11500 13151 11517
rect 13145 11497 13166 11500
rect 13163 11496 13166 11497
rect 13192 11496 13195 11522
rect 18545 11496 18548 11522
rect 18574 11516 18577 11522
rect 19604 11517 19633 11520
rect 19604 11516 19610 11517
rect 18574 11502 19610 11516
rect 18574 11496 18577 11502
rect 19604 11500 19610 11502
rect 19627 11500 19633 11517
rect 19604 11497 19633 11500
rect 9676 11468 10242 11482
rect 10311 11462 10314 11488
rect 10340 11462 10343 11488
rect 16107 11462 16110 11488
rect 16136 11482 16139 11488
rect 16338 11483 16367 11486
rect 16338 11482 16344 11483
rect 16136 11468 16344 11482
rect 16136 11462 16139 11468
rect 16338 11466 16344 11468
rect 16361 11466 16367 11483
rect 16338 11463 16367 11466
rect 3036 11400 29992 11448
rect 7597 11360 7600 11386
rect 7626 11380 7629 11386
rect 9667 11380 9670 11386
rect 7626 11366 9670 11380
rect 7626 11360 7629 11366
rect 9667 11360 9670 11366
rect 9696 11360 9699 11386
rect 21513 11381 21542 11384
rect 21513 11364 21519 11381
rect 21536 11380 21542 11381
rect 21673 11380 21676 11386
rect 21536 11366 21676 11380
rect 21536 11364 21542 11366
rect 21513 11361 21542 11364
rect 21673 11360 21676 11366
rect 21702 11360 21705 11386
rect 24433 11360 24436 11386
rect 24462 11360 24465 11386
rect 4745 11350 4748 11352
rect 4727 11347 4748 11350
rect 4727 11330 4733 11347
rect 4727 11327 4748 11330
rect 4745 11326 4748 11327
rect 4774 11326 4777 11352
rect 5757 11326 5760 11352
rect 5786 11346 5789 11352
rect 6171 11346 6174 11352
rect 5786 11332 6174 11346
rect 5786 11326 5789 11332
rect 6171 11326 6174 11332
rect 6200 11346 6203 11352
rect 6746 11347 6775 11350
rect 6746 11346 6752 11347
rect 6200 11332 6752 11346
rect 6200 11326 6203 11332
rect 6746 11330 6752 11332
rect 6769 11330 6775 11347
rect 6746 11327 6775 11330
rect 6797 11347 6826 11350
rect 6797 11330 6803 11347
rect 6820 11346 6826 11347
rect 6861 11346 6864 11352
rect 6820 11332 6864 11346
rect 6820 11330 6826 11332
rect 6797 11327 6826 11330
rect 6861 11326 6864 11332
rect 6890 11326 6893 11352
rect 17488 11347 17517 11350
rect 17488 11346 17494 11347
rect 16208 11332 17494 11346
rect 4515 11292 4518 11318
rect 4544 11292 4547 11318
rect 4677 11313 4706 11316
rect 4677 11296 4683 11313
rect 4700 11312 4706 11313
rect 6401 11312 6404 11318
rect 4700 11298 6404 11312
rect 4700 11296 4706 11298
rect 4677 11293 4706 11296
rect 6401 11292 6404 11298
rect 6430 11292 6433 11318
rect 16153 11292 16156 11318
rect 16182 11312 16185 11318
rect 16208 11316 16222 11332
rect 17488 11330 17494 11332
rect 17511 11330 17517 11347
rect 18591 11346 18594 11352
rect 17488 11327 17517 11330
rect 18462 11332 18594 11346
rect 16200 11313 16229 11316
rect 16200 11312 16206 11313
rect 16182 11298 16206 11312
rect 16182 11292 16185 11298
rect 16200 11296 16206 11298
rect 16223 11296 16229 11313
rect 16200 11293 16229 11296
rect 16292 11313 16321 11316
rect 16292 11296 16298 11313
rect 16315 11312 16321 11313
rect 16567 11312 16570 11318
rect 16315 11298 16570 11312
rect 16315 11296 16321 11298
rect 16292 11293 16321 11296
rect 16567 11292 16570 11298
rect 16596 11312 16599 11318
rect 17119 11312 17122 11318
rect 16596 11298 17122 11312
rect 16596 11292 16599 11298
rect 17119 11292 17122 11298
rect 17148 11292 17151 11318
rect 17441 11292 17444 11318
rect 17470 11292 17473 11318
rect 17533 11292 17536 11318
rect 17562 11312 17565 11318
rect 18407 11312 18410 11318
rect 17562 11298 18410 11312
rect 17562 11292 17565 11298
rect 18407 11292 18410 11298
rect 18436 11292 18439 11318
rect 18462 11316 18476 11332
rect 18591 11326 18594 11332
rect 18620 11326 18623 11352
rect 20707 11350 20710 11352
rect 20689 11347 20710 11350
rect 20689 11330 20695 11347
rect 20689 11327 20710 11330
rect 20707 11326 20710 11327
rect 20736 11326 20739 11352
rect 28343 11350 28346 11352
rect 28325 11347 28346 11350
rect 28325 11330 28331 11347
rect 28372 11346 28375 11352
rect 29149 11347 29178 11350
rect 28372 11332 28458 11346
rect 28325 11327 28346 11330
rect 28343 11326 28346 11327
rect 28372 11326 28375 11332
rect 18454 11313 18483 11316
rect 18454 11296 18460 11313
rect 18477 11296 18483 11313
rect 18454 11293 18483 11296
rect 18545 11292 18548 11318
rect 18574 11292 18577 11318
rect 20109 11292 20112 11318
rect 20138 11312 20141 11318
rect 20633 11313 20662 11316
rect 20633 11312 20639 11313
rect 20138 11298 20639 11312
rect 20138 11292 20141 11298
rect 20633 11296 20639 11298
rect 20656 11296 20662 11313
rect 20633 11293 20662 11296
rect 24295 11292 24298 11318
rect 24324 11312 24327 11318
rect 24342 11313 24371 11316
rect 24342 11312 24348 11313
rect 24324 11298 24348 11312
rect 24324 11292 24327 11298
rect 24342 11296 24348 11298
rect 24365 11296 24371 11313
rect 24342 11293 24371 11296
rect 24480 11313 24509 11316
rect 24480 11296 24486 11313
rect 24503 11296 24509 11313
rect 24480 11293 24509 11296
rect 5619 11258 5622 11284
rect 5648 11278 5651 11284
rect 5895 11278 5898 11284
rect 5648 11264 5898 11278
rect 5648 11258 5651 11264
rect 5895 11258 5898 11264
rect 5924 11278 5927 11284
rect 6586 11279 6615 11282
rect 6586 11278 6592 11279
rect 5924 11264 6592 11278
rect 5924 11258 5927 11264
rect 6586 11262 6592 11264
rect 6609 11262 6615 11279
rect 6586 11259 6615 11262
rect 7551 11258 7554 11284
rect 7580 11278 7583 11284
rect 7621 11279 7650 11282
rect 7621 11278 7627 11279
rect 7580 11264 7627 11278
rect 7580 11258 7583 11264
rect 7621 11262 7627 11264
rect 7644 11262 7650 11279
rect 7621 11259 7650 11262
rect 17073 11258 17076 11284
rect 17102 11258 17105 11284
rect 17211 11258 17214 11284
rect 17240 11258 17243 11284
rect 16062 11245 16091 11248
rect 16062 11228 16068 11245
rect 16085 11244 16091 11245
rect 16245 11244 16248 11250
rect 16085 11230 16248 11244
rect 16085 11228 16091 11230
rect 16062 11225 16091 11228
rect 16245 11224 16248 11230
rect 16274 11244 16277 11250
rect 17166 11245 17195 11248
rect 17166 11244 17172 11245
rect 16274 11230 17172 11244
rect 16274 11224 16277 11230
rect 17166 11228 17172 11230
rect 17189 11228 17195 11245
rect 18554 11244 18568 11292
rect 20155 11258 20158 11284
rect 20184 11278 20187 11284
rect 20478 11279 20507 11282
rect 20478 11278 20484 11279
rect 20184 11264 20484 11278
rect 20184 11258 20187 11264
rect 20478 11262 20484 11264
rect 20501 11262 20507 11279
rect 24488 11278 24502 11293
rect 24571 11292 24574 11318
rect 24600 11292 24603 11318
rect 28275 11313 28304 11316
rect 28275 11296 28281 11313
rect 28298 11312 28304 11313
rect 28389 11312 28392 11318
rect 28298 11298 28392 11312
rect 28298 11296 28304 11298
rect 28275 11293 28304 11296
rect 28389 11292 28392 11298
rect 28418 11292 28421 11318
rect 28444 11312 28458 11332
rect 29149 11330 29155 11347
rect 29172 11346 29178 11347
rect 29172 11332 29516 11346
rect 29172 11330 29178 11332
rect 29149 11327 29178 11330
rect 28665 11312 28668 11318
rect 28444 11298 28668 11312
rect 28665 11292 28668 11298
rect 28694 11292 28697 11318
rect 28711 11292 28714 11318
rect 28740 11312 28743 11318
rect 28849 11312 28852 11318
rect 28740 11298 28852 11312
rect 28740 11292 28743 11298
rect 28849 11292 28852 11298
rect 28878 11312 28881 11318
rect 29502 11316 29516 11332
rect 29402 11313 29431 11316
rect 29402 11312 29408 11313
rect 28878 11298 29408 11312
rect 28878 11292 28881 11298
rect 29402 11296 29408 11298
rect 29425 11296 29431 11313
rect 29402 11293 29431 11296
rect 29494 11313 29523 11316
rect 29494 11296 29500 11313
rect 29517 11296 29523 11313
rect 29494 11293 29523 11296
rect 24755 11278 24758 11284
rect 24488 11264 24758 11278
rect 20478 11259 20507 11262
rect 17166 11225 17195 11228
rect 17220 11230 18568 11244
rect 5527 11190 5530 11216
rect 5556 11214 5559 11216
rect 5556 11211 5580 11214
rect 5556 11194 5557 11211
rect 5574 11194 5580 11211
rect 5556 11191 5580 11194
rect 5556 11190 5559 11191
rect 16199 11190 16202 11216
rect 16228 11190 16231 11216
rect 16337 11190 16340 11216
rect 16366 11210 16369 11216
rect 17220 11210 17234 11230
rect 16366 11196 17234 11210
rect 18500 11211 18529 11214
rect 16366 11190 16369 11196
rect 18500 11194 18506 11211
rect 18523 11210 18529 11211
rect 18591 11210 18594 11216
rect 18523 11196 18594 11210
rect 18523 11194 18529 11196
rect 18500 11191 18529 11194
rect 18591 11190 18594 11196
rect 18620 11190 18623 11216
rect 20486 11210 20500 11259
rect 24755 11258 24758 11264
rect 24784 11258 24787 11284
rect 28113 11258 28116 11284
rect 28142 11258 28145 11284
rect 21167 11210 21170 11216
rect 20486 11196 21170 11210
rect 21167 11190 21170 11196
rect 21196 11190 21199 11216
rect 29447 11190 29450 11216
rect 29476 11190 29479 11216
rect 3036 11128 29992 11176
rect 18454 11109 18483 11112
rect 18454 11092 18460 11109
rect 18477 11108 18483 11109
rect 18729 11108 18732 11114
rect 18477 11094 18732 11108
rect 18477 11092 18483 11094
rect 18454 11089 18483 11092
rect 18729 11088 18732 11094
rect 18758 11088 18761 11114
rect 24571 11088 24574 11114
rect 24600 11108 24603 11114
rect 29079 11108 29082 11114
rect 24600 11094 29082 11108
rect 24600 11088 24603 11094
rect 29079 11088 29082 11094
rect 29108 11088 29111 11114
rect 6655 11075 6684 11078
rect 6655 11058 6661 11075
rect 6678 11074 6684 11075
rect 7459 11074 7462 11080
rect 6678 11060 7462 11074
rect 6678 11058 6684 11060
rect 6655 11055 6684 11058
rect 7459 11054 7462 11060
rect 7488 11054 7491 11080
rect 16936 11075 16965 11078
rect 16936 11058 16942 11075
rect 16959 11074 16965 11075
rect 17027 11074 17030 11080
rect 16959 11060 17030 11074
rect 16959 11058 16965 11060
rect 16936 11055 16965 11058
rect 17027 11054 17030 11060
rect 17056 11054 17059 11080
rect 17119 11054 17122 11080
rect 17148 11074 17151 11080
rect 17148 11060 17280 11074
rect 17148 11054 17151 11060
rect 5343 11020 5346 11046
rect 5372 11020 5375 11046
rect 11829 11020 11832 11046
rect 11858 11044 11861 11046
rect 11858 11041 11882 11044
rect 11858 11024 11859 11041
rect 11876 11024 11882 11041
rect 11858 11021 11882 11024
rect 11858 11020 11861 11021
rect 13945 11020 13948 11046
rect 13974 11020 13977 11046
rect 16337 11020 16340 11046
rect 16366 11020 16369 11046
rect 17211 11020 17214 11046
rect 17240 11020 17243 11046
rect 5252 11007 5281 11010
rect 5252 10990 5258 11007
rect 5275 11006 5281 11007
rect 5527 11006 5530 11012
rect 5275 10992 5530 11006
rect 5275 10990 5281 10992
rect 5252 10987 5281 10990
rect 5527 10986 5530 10992
rect 5556 10986 5559 11012
rect 5619 10986 5622 11012
rect 5648 10986 5651 11012
rect 5757 10986 5760 11012
rect 5786 11010 5789 11012
rect 5786 11007 5804 11010
rect 5798 10990 5804 11007
rect 6907 11006 6910 11012
rect 5786 10987 5804 10990
rect 5950 10992 6910 11006
rect 5786 10986 5789 10987
rect 5831 10973 5860 10976
rect 5831 10956 5837 10973
rect 5854 10972 5860 10973
rect 5950 10972 5964 10992
rect 6907 10986 6910 10992
rect 6936 10986 6939 11012
rect 10035 10986 10038 11012
rect 10064 11006 10067 11012
rect 10818 11007 10847 11010
rect 10818 11006 10824 11007
rect 10064 10992 10824 11006
rect 10064 10986 10067 10992
rect 10818 10990 10824 10992
rect 10841 11006 10847 11007
rect 10863 11006 10866 11012
rect 10841 10992 10866 11006
rect 10841 10990 10847 10992
rect 10818 10987 10847 10990
rect 10863 10986 10866 10992
rect 10892 10986 10895 11012
rect 10979 11007 11008 11010
rect 10979 10990 10985 11007
rect 11002 11006 11008 11007
rect 11093 11006 11096 11012
rect 11002 10992 11096 11006
rect 11002 10990 11008 10992
rect 10979 10987 11008 10990
rect 11093 10986 11096 10992
rect 11122 10986 11125 11012
rect 12611 10986 12614 11012
rect 12640 11006 12643 11012
rect 14497 11006 14500 11012
rect 12640 10992 14500 11006
rect 12640 10986 12643 10992
rect 14497 10986 14500 10992
rect 14526 10986 14529 11012
rect 16153 10986 16156 11012
rect 16182 11006 16185 11012
rect 16200 11007 16229 11010
rect 16200 11006 16206 11007
rect 16182 10992 16206 11006
rect 16182 10986 16185 10992
rect 16200 10990 16206 10992
rect 16223 10990 16229 11007
rect 16200 10987 16229 10990
rect 16245 10986 16248 11012
rect 16274 10986 16277 11012
rect 16383 10986 16386 11012
rect 16412 11006 16415 11012
rect 16890 11007 16919 11010
rect 16890 11006 16896 11007
rect 16412 10992 16896 11006
rect 16412 10986 16415 10992
rect 16890 10990 16896 10992
rect 16913 10990 16919 11007
rect 16890 10987 16919 10990
rect 11047 10976 11050 10978
rect 5854 10958 5964 10972
rect 11029 10973 11050 10976
rect 5854 10956 5860 10958
rect 5831 10953 5860 10956
rect 11029 10956 11035 10973
rect 11029 10953 11050 10956
rect 11047 10952 11050 10953
rect 11076 10952 11079 10978
rect 16898 10972 16912 10987
rect 17165 10986 17168 11012
rect 17194 10986 17197 11012
rect 17266 11006 17280 11060
rect 21167 11020 21170 11046
rect 21196 11040 21199 11046
rect 21214 11041 21243 11044
rect 21214 11040 21220 11041
rect 21196 11026 21220 11040
rect 21196 11020 21199 11026
rect 21214 11024 21220 11026
rect 21237 11024 21243 11041
rect 21214 11021 21243 11024
rect 22087 11020 22090 11046
rect 22116 11040 22119 11046
rect 22502 11041 22531 11044
rect 22502 11040 22508 11041
rect 22116 11026 22508 11040
rect 22116 11020 22119 11026
rect 22502 11024 22508 11026
rect 22525 11024 22531 11041
rect 22502 11021 22531 11024
rect 22915 11020 22918 11046
rect 22944 11040 22947 11046
rect 26687 11040 26690 11046
rect 22944 11026 26690 11040
rect 22944 11020 22947 11026
rect 26687 11020 26690 11026
rect 26716 11020 26719 11046
rect 17901 11006 17904 11012
rect 17266 10992 17904 11006
rect 17901 10986 17904 10992
rect 17930 11006 17933 11012
rect 18454 11007 18483 11010
rect 18454 11006 18460 11007
rect 17930 10992 18460 11006
rect 17930 10986 17933 10992
rect 18454 10990 18460 10992
rect 18477 10990 18483 11007
rect 18454 10987 18483 10990
rect 18591 10986 18594 11012
rect 18620 10986 18623 11012
rect 22685 10986 22688 11012
rect 22714 11010 22717 11012
rect 22714 11006 22718 11010
rect 22714 10992 22736 11006
rect 22714 10987 22718 10992
rect 22714 10986 22717 10987
rect 23145 10986 23148 11012
rect 23174 10986 23177 11012
rect 23237 10986 23240 11012
rect 23266 10986 23269 11012
rect 23973 10986 23976 11012
rect 24002 10986 24005 11012
rect 24066 11007 24095 11010
rect 24066 10990 24072 11007
rect 24089 10990 24095 11007
rect 24066 10987 24095 10990
rect 17257 10972 17260 10978
rect 16898 10958 17260 10972
rect 17257 10952 17260 10958
rect 17286 10952 17289 10978
rect 18315 10952 18318 10978
rect 18344 10972 18347 10978
rect 18546 10973 18575 10976
rect 18546 10972 18552 10973
rect 18344 10958 18552 10972
rect 18344 10952 18347 10958
rect 18546 10956 18552 10958
rect 18569 10956 18575 10973
rect 18546 10953 18575 10956
rect 21213 10952 21216 10978
rect 21242 10972 21245 10978
rect 21443 10976 21446 10978
rect 21374 10973 21403 10976
rect 21374 10972 21380 10973
rect 21242 10958 21380 10972
rect 21242 10952 21245 10958
rect 21374 10956 21380 10958
rect 21397 10956 21403 10973
rect 21374 10953 21403 10956
rect 21425 10973 21446 10976
rect 21425 10956 21431 10973
rect 21425 10953 21446 10956
rect 21443 10952 21446 10953
rect 21472 10952 21475 10978
rect 22249 10973 22278 10976
rect 22249 10956 22255 10973
rect 22272 10972 22278 10973
rect 22502 10973 22531 10976
rect 22502 10972 22508 10973
rect 22272 10958 22508 10972
rect 22272 10956 22278 10958
rect 22249 10953 22278 10956
rect 22502 10956 22508 10958
rect 22525 10956 22531 10973
rect 22502 10953 22531 10956
rect 22593 10952 22596 10978
rect 22622 10952 22625 10978
rect 22639 10952 22642 10978
rect 22668 10952 22671 10978
rect 23007 10952 23010 10978
rect 23036 10972 23039 10978
rect 24074 10972 24088 10987
rect 23036 10958 24088 10972
rect 23036 10952 23039 10958
rect 5022 10939 5051 10942
rect 5022 10922 5028 10939
rect 5045 10938 5051 10939
rect 5113 10938 5116 10944
rect 5045 10924 5116 10938
rect 5045 10922 5051 10924
rect 5022 10919 5051 10922
rect 5113 10918 5116 10924
rect 5142 10918 5145 10944
rect 5205 10918 5208 10944
rect 5234 10918 5237 10944
rect 13669 10918 13672 10944
rect 13698 10918 13701 10944
rect 13853 10918 13856 10944
rect 13882 10918 13885 10944
rect 13899 10918 13902 10944
rect 13928 10918 13931 10944
rect 15877 10918 15880 10944
rect 15906 10938 15909 10944
rect 16108 10939 16137 10942
rect 16108 10938 16114 10939
rect 15906 10924 16114 10938
rect 15906 10918 15909 10924
rect 16108 10922 16114 10924
rect 16131 10922 16137 10939
rect 16108 10919 16137 10922
rect 23191 10918 23194 10944
rect 23220 10918 23223 10944
rect 24019 10918 24022 10944
rect 24048 10918 24051 10944
rect 3036 10856 29992 10904
rect 13417 10837 13446 10840
rect 11036 10822 12220 10836
rect 4745 10782 4748 10808
rect 4774 10802 4777 10808
rect 10243 10803 10272 10806
rect 10243 10802 10249 10803
rect 4774 10788 10249 10802
rect 4774 10782 4777 10788
rect 10243 10786 10249 10788
rect 10266 10802 10272 10803
rect 10266 10788 10380 10802
rect 10266 10786 10272 10788
rect 10243 10783 10272 10786
rect 10035 10748 10038 10774
rect 10064 10748 10067 10774
rect 10197 10769 10226 10772
rect 10197 10752 10203 10769
rect 10220 10768 10226 10769
rect 10311 10768 10314 10774
rect 10220 10754 10314 10768
rect 10220 10752 10226 10754
rect 10197 10749 10226 10752
rect 10311 10748 10314 10754
rect 10340 10748 10343 10774
rect 10366 10768 10380 10788
rect 11036 10768 11050 10822
rect 11071 10803 11100 10806
rect 11071 10786 11077 10803
rect 11094 10802 11100 10803
rect 11094 10788 12174 10802
rect 11094 10786 11100 10788
rect 11071 10783 11100 10786
rect 12160 10772 12174 10788
rect 10366 10754 11050 10768
rect 11830 10769 11859 10772
rect 11830 10752 11836 10769
rect 11853 10768 11859 10769
rect 12152 10769 12181 10772
rect 11853 10754 11990 10768
rect 11853 10752 11859 10754
rect 11830 10749 11859 10752
rect 11875 10714 11878 10740
rect 11904 10734 11907 10740
rect 11922 10735 11951 10738
rect 11922 10734 11928 10735
rect 11904 10720 11928 10734
rect 11904 10714 11907 10720
rect 11922 10718 11928 10720
rect 11945 10718 11951 10735
rect 11922 10715 11951 10718
rect 11976 10700 11990 10754
rect 12152 10752 12158 10769
rect 12175 10752 12181 10769
rect 12206 10768 12220 10822
rect 13417 10820 13423 10837
rect 13440 10836 13446 10837
rect 13899 10836 13902 10842
rect 13440 10822 13902 10836
rect 13440 10820 13446 10822
rect 13417 10817 13446 10820
rect 13899 10816 13902 10822
rect 13928 10816 13931 10842
rect 15739 10816 15742 10842
rect 15768 10836 15771 10842
rect 15786 10837 15815 10840
rect 15786 10836 15792 10837
rect 15768 10822 15792 10836
rect 15768 10816 15771 10822
rect 15786 10820 15792 10822
rect 15809 10820 15815 10837
rect 15786 10817 15815 10820
rect 16521 10816 16524 10842
rect 16550 10836 16553 10842
rect 20339 10836 20342 10842
rect 16550 10822 20342 10836
rect 16550 10816 16553 10822
rect 20339 10816 20342 10822
rect 20368 10816 20371 10842
rect 22111 10837 22140 10840
rect 22111 10820 22117 10837
rect 22134 10836 22140 10837
rect 22639 10836 22642 10842
rect 22134 10822 22642 10836
rect 22134 10820 22140 10822
rect 22111 10817 22140 10820
rect 22639 10816 22642 10822
rect 22668 10816 22671 10842
rect 22962 10837 22991 10840
rect 22962 10820 22968 10837
rect 22985 10836 22991 10837
rect 23237 10836 23240 10842
rect 22985 10822 23240 10836
rect 22985 10820 22991 10822
rect 22962 10817 22991 10820
rect 23237 10816 23240 10822
rect 23266 10816 23269 10842
rect 23513 10816 23516 10842
rect 23542 10836 23545 10842
rect 23542 10822 24364 10836
rect 23542 10816 23545 10822
rect 12427 10782 12430 10808
rect 12456 10802 12459 10808
rect 12611 10806 12614 10808
rect 12542 10803 12571 10806
rect 12542 10802 12548 10803
rect 12456 10788 12548 10802
rect 12456 10782 12459 10788
rect 12542 10786 12548 10788
rect 12565 10786 12571 10803
rect 12542 10783 12571 10786
rect 12593 10803 12614 10806
rect 12593 10786 12599 10803
rect 12593 10783 12614 10786
rect 12600 10768 12614 10783
rect 12640 10782 12643 10808
rect 14497 10782 14500 10808
rect 14526 10802 14529 10808
rect 14663 10803 14692 10806
rect 14663 10802 14669 10803
rect 14526 10788 14669 10802
rect 14526 10782 14529 10788
rect 14663 10786 14669 10788
rect 14686 10802 14692 10803
rect 15487 10803 15516 10806
rect 14686 10788 14796 10802
rect 14686 10786 14692 10788
rect 14663 10783 14692 10786
rect 12206 10754 12614 10768
rect 14613 10769 14642 10772
rect 12152 10749 12181 10752
rect 14613 10752 14619 10769
rect 14636 10768 14642 10769
rect 14727 10768 14730 10774
rect 14636 10754 14730 10768
rect 14636 10752 14642 10754
rect 14613 10749 14642 10752
rect 14727 10748 14730 10754
rect 14756 10748 14759 10774
rect 14782 10768 14796 10788
rect 15487 10786 15493 10803
rect 15510 10802 15516 10803
rect 15510 10788 16222 10802
rect 15510 10786 15516 10788
rect 15487 10783 15516 10786
rect 15141 10768 15144 10774
rect 14782 10754 15144 10768
rect 15141 10748 15144 10754
rect 15170 10748 15173 10774
rect 16208 10772 16222 10788
rect 18278 10788 19396 10802
rect 18278 10772 18292 10788
rect 15786 10769 15815 10772
rect 15786 10768 15792 10769
rect 15334 10754 15792 10768
rect 12381 10714 12384 10740
rect 12410 10714 12413 10740
rect 14037 10714 14040 10740
rect 14066 10734 14069 10740
rect 14452 10735 14481 10738
rect 14452 10734 14458 10735
rect 14066 10720 14458 10734
rect 14066 10714 14069 10720
rect 14452 10718 14458 10720
rect 14475 10718 14481 10735
rect 14452 10715 14481 10718
rect 11976 10686 12082 10700
rect 5343 10646 5346 10672
rect 5372 10666 5375 10672
rect 10679 10666 10682 10672
rect 5372 10652 10682 10666
rect 5372 10646 5375 10652
rect 10679 10646 10682 10652
rect 10708 10646 10711 10672
rect 12068 10666 12082 10686
rect 15334 10666 15348 10754
rect 15786 10752 15792 10754
rect 15809 10768 15815 10769
rect 16200 10769 16229 10772
rect 15809 10754 15877 10768
rect 15809 10752 15815 10754
rect 15786 10749 15815 10752
rect 15863 10734 15877 10754
rect 16200 10752 16206 10769
rect 16223 10752 16229 10769
rect 16200 10749 16229 10752
rect 18270 10769 18299 10772
rect 18270 10752 18276 10769
rect 18293 10752 18299 10769
rect 18270 10749 18299 10752
rect 18729 10748 18732 10774
rect 18758 10768 18761 10774
rect 18812 10769 18841 10772
rect 18812 10768 18818 10769
rect 18758 10754 18818 10768
rect 18758 10748 18761 10754
rect 18812 10752 18818 10754
rect 18835 10752 18841 10769
rect 18812 10749 18841 10752
rect 17533 10734 17536 10740
rect 15863 10720 17536 10734
rect 17533 10714 17536 10720
rect 17562 10714 17565 10740
rect 18315 10714 18318 10740
rect 18344 10714 18347 10740
rect 18684 10735 18713 10738
rect 18684 10718 18690 10735
rect 18707 10718 18713 10735
rect 18684 10715 18713 10718
rect 12068 10652 15348 10666
rect 18408 10667 18437 10670
rect 18408 10650 18414 10667
rect 18431 10666 18437 10667
rect 18637 10666 18640 10672
rect 18431 10652 18640 10666
rect 18431 10650 18437 10652
rect 18408 10647 18437 10650
rect 18637 10646 18640 10652
rect 18666 10646 18669 10672
rect 18692 10666 18706 10715
rect 19382 10704 19396 10788
rect 19925 10782 19928 10808
rect 19954 10802 19957 10808
rect 20202 10803 20231 10806
rect 20202 10802 20208 10803
rect 19954 10788 20208 10802
rect 19954 10782 19957 10788
rect 20202 10786 20208 10788
rect 20225 10786 20231 10803
rect 20202 10783 20231 10786
rect 20891 10782 20894 10808
rect 20920 10802 20923 10808
rect 21275 10803 21304 10806
rect 21275 10802 21281 10803
rect 20920 10788 21281 10802
rect 20920 10782 20923 10788
rect 21275 10786 21281 10788
rect 21298 10802 21304 10803
rect 21351 10802 21354 10808
rect 21298 10788 21354 10802
rect 21298 10786 21304 10788
rect 21275 10783 21304 10786
rect 21351 10782 21354 10788
rect 21380 10782 21383 10808
rect 23191 10782 23194 10808
rect 23220 10802 23223 10808
rect 23361 10803 23390 10806
rect 23361 10802 23367 10803
rect 23220 10788 23367 10802
rect 23220 10782 23223 10788
rect 23361 10786 23367 10788
rect 23384 10786 23390 10803
rect 23361 10783 23390 10786
rect 24019 10782 24022 10808
rect 24048 10802 24051 10808
rect 24281 10803 24310 10806
rect 24281 10802 24287 10803
rect 24048 10788 24287 10802
rect 24048 10782 24051 10788
rect 24281 10786 24287 10788
rect 24304 10786 24310 10803
rect 24350 10802 24364 10822
rect 26825 10816 26828 10842
rect 26854 10816 26857 10842
rect 29079 10816 29082 10842
rect 29108 10816 29111 10842
rect 25583 10806 25586 10808
rect 25565 10803 25586 10806
rect 25565 10802 25571 10803
rect 24350 10788 25571 10802
rect 24281 10783 24310 10786
rect 25565 10786 25571 10788
rect 25565 10783 25586 10786
rect 25583 10782 25586 10783
rect 25612 10782 25615 10808
rect 29126 10803 29155 10806
rect 29126 10786 29132 10803
rect 29149 10802 29155 10803
rect 29493 10802 29496 10808
rect 29149 10788 29496 10802
rect 29149 10786 29155 10788
rect 29126 10783 29155 10786
rect 29493 10782 29496 10788
rect 29522 10782 29525 10808
rect 20293 10748 20296 10774
rect 20322 10748 20325 10774
rect 20340 10769 20369 10772
rect 20340 10752 20346 10769
rect 20363 10768 20369 10769
rect 20431 10768 20434 10774
rect 20363 10754 20434 10768
rect 20363 10752 20369 10754
rect 20340 10749 20369 10752
rect 20431 10748 20434 10754
rect 20460 10748 20463 10774
rect 21213 10768 21216 10774
rect 21242 10772 21245 10774
rect 21242 10769 21260 10772
rect 20578 10754 21216 10768
rect 20109 10714 20112 10740
rect 20138 10734 20141 10740
rect 20578 10734 20592 10754
rect 21213 10748 21216 10754
rect 21254 10752 21260 10769
rect 21242 10749 21260 10752
rect 21242 10748 21245 10749
rect 22915 10748 22918 10774
rect 22944 10748 22947 10774
rect 23008 10769 23037 10772
rect 23008 10752 23014 10769
rect 23031 10768 23037 10769
rect 23099 10768 23102 10774
rect 23031 10754 23102 10768
rect 23031 10752 23037 10754
rect 23008 10749 23037 10752
rect 23099 10748 23102 10754
rect 23128 10748 23131 10774
rect 25515 10769 25544 10772
rect 23246 10754 23766 10768
rect 23246 10740 23260 10754
rect 20138 10720 20592 10734
rect 21076 10735 21105 10738
rect 20138 10714 20141 10720
rect 21076 10718 21082 10735
rect 21099 10718 21105 10735
rect 21076 10715 21105 10718
rect 19374 10701 19403 10704
rect 19374 10684 19380 10701
rect 19397 10700 19403 10701
rect 19925 10700 19928 10706
rect 19397 10686 19928 10700
rect 19397 10684 19403 10686
rect 19374 10681 19403 10684
rect 19925 10680 19928 10686
rect 19954 10680 19957 10706
rect 19327 10666 19330 10672
rect 18692 10652 19330 10666
rect 19327 10646 19330 10652
rect 19356 10666 19359 10672
rect 20155 10666 20158 10672
rect 19356 10652 20158 10666
rect 19356 10646 19359 10652
rect 20155 10646 20158 10652
rect 20184 10646 20187 10672
rect 20202 10667 20231 10670
rect 20202 10650 20208 10667
rect 20225 10666 20231 10667
rect 20615 10666 20618 10672
rect 20225 10652 20618 10666
rect 20225 10650 20231 10652
rect 20202 10647 20231 10650
rect 20615 10646 20618 10652
rect 20644 10646 20647 10672
rect 21084 10666 21098 10715
rect 23237 10714 23240 10740
rect 23266 10714 23269 10740
rect 23752 10734 23766 10754
rect 25515 10752 25521 10769
rect 25538 10768 25544 10769
rect 25675 10768 25678 10774
rect 25538 10754 25678 10768
rect 25538 10752 25544 10754
rect 25515 10749 25544 10752
rect 25675 10748 25678 10754
rect 25704 10748 25707 10774
rect 26688 10769 26717 10772
rect 26688 10752 26694 10769
rect 26711 10768 26717 10769
rect 27009 10768 27012 10774
rect 26711 10754 27012 10768
rect 26711 10752 26717 10754
rect 26688 10749 26717 10752
rect 27009 10748 27012 10754
rect 27038 10748 27041 10774
rect 28941 10748 28944 10774
rect 28970 10768 28973 10774
rect 29034 10769 29063 10772
rect 29034 10768 29040 10769
rect 28970 10754 29040 10768
rect 28970 10748 28973 10754
rect 29034 10752 29040 10754
rect 29057 10752 29063 10769
rect 29034 10749 29063 10752
rect 29172 10769 29201 10772
rect 29172 10752 29178 10769
rect 29195 10768 29201 10769
rect 29447 10768 29450 10774
rect 29195 10754 29450 10768
rect 29195 10752 29201 10754
rect 29172 10749 29201 10752
rect 29447 10748 29450 10754
rect 29476 10748 29479 10774
rect 24158 10735 24187 10738
rect 24158 10734 24164 10735
rect 23752 10720 24164 10734
rect 24158 10718 24164 10720
rect 24181 10718 24187 10735
rect 24158 10715 24187 10718
rect 21167 10666 21170 10672
rect 21084 10652 21170 10666
rect 21167 10646 21170 10652
rect 21196 10666 21199 10672
rect 23237 10666 23240 10672
rect 21196 10652 23240 10666
rect 21196 10646 21199 10652
rect 23237 10646 23240 10652
rect 23266 10646 23269 10672
rect 23559 10646 23562 10672
rect 23588 10666 23591 10672
rect 23928 10667 23957 10670
rect 23928 10666 23934 10667
rect 23588 10652 23934 10666
rect 23588 10646 23591 10652
rect 23928 10650 23934 10652
rect 23951 10650 23957 10667
rect 24166 10666 24180 10715
rect 24663 10714 24666 10740
rect 24692 10734 24695 10740
rect 24801 10734 24804 10740
rect 24692 10720 24804 10734
rect 24692 10714 24695 10720
rect 24801 10714 24804 10720
rect 24830 10714 24833 10740
rect 25353 10734 25356 10740
rect 24856 10720 25356 10734
rect 24856 10700 24870 10720
rect 25353 10714 25356 10720
rect 25382 10714 25385 10740
rect 26227 10714 26230 10740
rect 26256 10734 26259 10740
rect 26826 10735 26855 10738
rect 26826 10734 26832 10735
rect 26256 10720 26832 10734
rect 26256 10714 26259 10720
rect 26826 10718 26832 10720
rect 26849 10718 26855 10735
rect 26826 10715 26855 10718
rect 24626 10686 24870 10700
rect 24626 10672 24640 10686
rect 24617 10666 24620 10672
rect 24166 10652 24620 10666
rect 23928 10647 23957 10650
rect 24617 10646 24620 10652
rect 24646 10646 24649 10672
rect 24848 10667 24877 10670
rect 24848 10650 24854 10667
rect 24871 10666 24877 10667
rect 24893 10666 24896 10672
rect 24871 10652 24896 10666
rect 24871 10650 24877 10652
rect 24848 10647 24877 10650
rect 24893 10646 24896 10652
rect 24922 10666 24925 10672
rect 25675 10666 25678 10672
rect 24922 10652 25678 10666
rect 24922 10646 24925 10652
rect 25675 10646 25678 10652
rect 25704 10646 25707 10672
rect 26273 10646 26276 10672
rect 26302 10666 26305 10672
rect 26389 10667 26418 10670
rect 26389 10666 26395 10667
rect 26302 10652 26395 10666
rect 26302 10646 26305 10652
rect 26389 10650 26395 10652
rect 26412 10650 26418 10667
rect 26389 10647 26418 10650
rect 26733 10646 26736 10672
rect 26762 10646 26765 10672
rect 3036 10584 29992 10632
rect 5619 10564 5622 10570
rect 4984 10550 5622 10564
rect 4984 10500 4998 10550
rect 5619 10544 5622 10550
rect 5648 10544 5651 10570
rect 9253 10564 9256 10570
rect 8526 10550 9256 10564
rect 4976 10497 5005 10500
rect 4976 10480 4982 10497
rect 4999 10480 5005 10497
rect 4976 10477 5005 10480
rect 5113 10476 5116 10502
rect 5142 10476 5145 10502
rect 8426 10497 8455 10500
rect 8426 10480 8432 10497
rect 8449 10496 8455 10497
rect 8471 10496 8474 10502
rect 8449 10482 8474 10496
rect 8449 10480 8455 10482
rect 8426 10477 8455 10480
rect 8471 10476 8474 10482
rect 8500 10476 8503 10502
rect 5665 10442 5668 10468
rect 5694 10462 5697 10468
rect 7597 10462 7600 10468
rect 5694 10448 7600 10462
rect 5694 10442 5697 10448
rect 7597 10442 7600 10448
rect 7626 10442 7629 10468
rect 8333 10442 8336 10468
rect 8362 10442 8365 10468
rect 8526 10466 8540 10550
rect 9253 10544 9256 10550
rect 9282 10544 9285 10570
rect 10679 10544 10682 10570
rect 10708 10564 10711 10570
rect 13945 10564 13948 10570
rect 10708 10550 13948 10564
rect 10708 10544 10711 10550
rect 13945 10544 13948 10550
rect 13974 10544 13977 10570
rect 17166 10565 17195 10568
rect 17166 10548 17172 10565
rect 17189 10564 17195 10565
rect 17257 10564 17260 10570
rect 17189 10550 17260 10564
rect 17189 10548 17195 10550
rect 17166 10545 17195 10548
rect 17257 10544 17260 10550
rect 17286 10544 17289 10570
rect 18684 10565 18713 10568
rect 18684 10548 18690 10565
rect 18707 10564 18713 10565
rect 18729 10564 18732 10570
rect 18707 10550 18732 10564
rect 18707 10548 18713 10550
rect 18684 10545 18713 10548
rect 18729 10544 18732 10550
rect 18758 10544 18761 10570
rect 20293 10544 20296 10570
rect 20322 10564 20325 10570
rect 20409 10565 20438 10568
rect 20409 10564 20415 10565
rect 20322 10550 20415 10564
rect 20322 10544 20325 10550
rect 20409 10548 20415 10550
rect 20432 10548 20438 10565
rect 20409 10545 20438 10548
rect 23007 10544 23010 10570
rect 23036 10544 23039 10570
rect 23145 10544 23148 10570
rect 23174 10564 23177 10570
rect 23422 10565 23451 10568
rect 23422 10564 23428 10565
rect 23174 10550 23428 10564
rect 23174 10544 23177 10550
rect 23422 10548 23428 10550
rect 23445 10548 23451 10565
rect 23422 10545 23451 10548
rect 23973 10544 23976 10570
rect 24002 10564 24005 10570
rect 24066 10565 24095 10568
rect 24066 10564 24072 10565
rect 24002 10550 24072 10564
rect 24002 10544 24005 10550
rect 24066 10548 24072 10550
rect 24089 10548 24095 10565
rect 24066 10545 24095 10548
rect 24111 10544 24114 10570
rect 24140 10564 24143 10570
rect 24140 10544 24157 10564
rect 14773 10510 14776 10536
rect 14802 10510 14805 10536
rect 20339 10510 20342 10536
rect 20368 10530 20371 10536
rect 24143 10530 24157 10544
rect 24626 10550 25537 10564
rect 24626 10530 24640 10550
rect 20368 10516 23490 10530
rect 24143 10516 24640 10530
rect 20368 10510 20371 10516
rect 8748 10497 8777 10500
rect 8748 10480 8754 10497
rect 8771 10496 8777 10497
rect 9529 10496 9532 10502
rect 8771 10482 9532 10496
rect 8771 10480 8777 10482
rect 8748 10477 8777 10480
rect 9529 10476 9532 10482
rect 9558 10476 9561 10502
rect 13669 10476 13672 10502
rect 13698 10476 13701 10502
rect 13853 10476 13856 10502
rect 13882 10496 13885 10502
rect 13945 10496 13948 10502
rect 13882 10482 13948 10496
rect 13882 10476 13885 10482
rect 13945 10476 13948 10482
rect 13974 10496 13977 10502
rect 14544 10497 14573 10500
rect 14544 10496 14550 10497
rect 13974 10482 14550 10496
rect 13974 10476 13977 10482
rect 14544 10480 14550 10482
rect 14567 10480 14573 10497
rect 14544 10477 14573 10480
rect 16016 10497 16045 10500
rect 16016 10480 16022 10497
rect 16039 10496 16045 10497
rect 16199 10496 16202 10502
rect 16039 10482 16202 10496
rect 16039 10480 16045 10482
rect 16016 10477 16045 10480
rect 16199 10476 16202 10482
rect 16228 10476 16231 10502
rect 19327 10476 19330 10502
rect 19356 10496 19359 10502
rect 23476 10500 23490 10516
rect 19374 10497 19403 10500
rect 19374 10496 19380 10497
rect 19356 10482 19380 10496
rect 19356 10476 19359 10482
rect 19374 10480 19380 10482
rect 19397 10480 19403 10497
rect 19374 10477 19403 10480
rect 23468 10497 23497 10500
rect 23468 10480 23474 10497
rect 23491 10496 23497 10497
rect 24112 10497 24141 10500
rect 24112 10496 24118 10497
rect 23491 10482 24118 10496
rect 23491 10480 23497 10482
rect 23468 10477 23497 10480
rect 24112 10480 24118 10482
rect 24135 10480 24141 10497
rect 24112 10477 24141 10480
rect 24617 10476 24620 10502
rect 24646 10476 24649 10502
rect 8518 10463 8547 10466
rect 8518 10446 8524 10463
rect 8541 10446 8547 10463
rect 8518 10443 8547 10446
rect 12381 10442 12384 10468
rect 12410 10462 12413 10468
rect 13532 10463 13561 10466
rect 13532 10462 13538 10463
rect 12410 10448 13538 10462
rect 12410 10442 12413 10448
rect 13532 10446 13538 10448
rect 13555 10446 13561 10463
rect 13532 10443 13561 10446
rect 5988 10429 6017 10432
rect 5988 10412 5994 10429
rect 6011 10412 6017 10429
rect 5988 10409 6017 10412
rect 8886 10429 8915 10432
rect 8886 10412 8892 10429
rect 8909 10428 8915 10429
rect 9023 10428 9026 10434
rect 8909 10414 9026 10428
rect 8909 10412 8915 10414
rect 8886 10409 8915 10412
rect 5205 10374 5208 10400
rect 5234 10394 5237 10400
rect 5996 10394 6010 10409
rect 9023 10408 9026 10414
rect 9052 10408 9055 10434
rect 9575 10428 9578 10434
rect 9499 10414 9578 10428
rect 9575 10408 9578 10414
rect 9604 10408 9607 10434
rect 5234 10380 6010 10394
rect 5234 10374 5237 10380
rect 8379 10374 8382 10400
rect 8408 10374 8411 10400
rect 8472 10395 8501 10398
rect 8472 10378 8478 10395
rect 8495 10394 8501 10395
rect 8931 10394 8934 10400
rect 8495 10380 8934 10394
rect 8495 10378 8501 10380
rect 8472 10375 8501 10378
rect 8931 10374 8934 10380
rect 8960 10374 8963 10400
rect 9253 10374 9256 10400
rect 9282 10394 9285 10400
rect 9622 10395 9651 10398
rect 9622 10394 9628 10395
rect 9282 10380 9628 10394
rect 9282 10374 9285 10380
rect 9622 10378 9628 10380
rect 9645 10378 9651 10395
rect 13540 10394 13554 10443
rect 14405 10442 14408 10468
rect 14434 10462 14437 10468
rect 14912 10463 14941 10466
rect 14912 10462 14918 10463
rect 14434 10448 14918 10462
rect 14434 10442 14437 10448
rect 14912 10446 14918 10448
rect 14935 10462 14941 10463
rect 15785 10462 15788 10468
rect 14935 10448 15788 10462
rect 14935 10446 14941 10448
rect 14912 10443 14941 10446
rect 15785 10442 15788 10448
rect 15814 10442 15817 10468
rect 15878 10463 15907 10466
rect 15878 10446 15884 10463
rect 15901 10446 15907 10463
rect 15878 10443 15907 10446
rect 13899 10408 13902 10434
rect 13928 10408 13931 10434
rect 14313 10428 14316 10434
rect 14283 10414 14316 10428
rect 14313 10408 14316 10414
rect 14342 10408 14345 10434
rect 14589 10408 14592 10434
rect 14618 10428 14621 10434
rect 14774 10429 14803 10432
rect 14774 10428 14780 10429
rect 14618 10414 14780 10428
rect 14618 10408 14621 10414
rect 14774 10412 14780 10414
rect 14797 10412 14803 10429
rect 15886 10428 15900 10443
rect 17211 10442 17214 10468
rect 17240 10442 17243 10468
rect 17396 10463 17425 10466
rect 17396 10446 17402 10463
rect 17419 10446 17425 10463
rect 17396 10443 17425 10446
rect 15969 10428 15972 10434
rect 15886 10414 15972 10428
rect 14774 10409 14803 10412
rect 15969 10408 15972 10414
rect 15998 10408 16001 10434
rect 16245 10408 16248 10434
rect 16274 10408 16277 10434
rect 16521 10408 16524 10434
rect 16550 10408 16553 10434
rect 16890 10429 16919 10432
rect 16890 10412 16896 10429
rect 16913 10412 16919 10429
rect 17404 10428 17418 10443
rect 18637 10442 18640 10468
rect 18666 10442 18669 10468
rect 18683 10442 18686 10468
rect 18712 10462 18715 10468
rect 18730 10463 18759 10466
rect 18730 10462 18736 10463
rect 18712 10448 18736 10462
rect 18712 10442 18715 10448
rect 18730 10446 18736 10448
rect 18753 10446 18759 10463
rect 18730 10443 18759 10446
rect 19535 10463 19564 10466
rect 19535 10446 19541 10463
rect 19558 10462 19564 10463
rect 20109 10462 20112 10468
rect 19558 10448 20112 10462
rect 19558 10446 19564 10448
rect 19535 10443 19564 10446
rect 20109 10442 20112 10448
rect 20138 10442 20141 10468
rect 23008 10463 23037 10466
rect 23008 10462 23014 10463
rect 20693 10448 23014 10462
rect 16890 10409 16919 10412
rect 17128 10414 17418 10428
rect 19585 10429 19614 10432
rect 14037 10394 14040 10400
rect 13540 10380 14040 10394
rect 9622 10375 9651 10378
rect 14037 10374 14040 10380
rect 14066 10374 14069 10400
rect 14865 10374 14868 10400
rect 14894 10374 14897 10400
rect 16898 10394 16912 10409
rect 17128 10400 17142 10414
rect 19585 10412 19591 10429
rect 19608 10428 19614 10429
rect 19649 10428 19652 10434
rect 19608 10414 19652 10428
rect 19608 10412 19614 10414
rect 19585 10409 19614 10412
rect 19649 10408 19652 10414
rect 19678 10408 19681 10434
rect 17119 10394 17122 10400
rect 16898 10380 17122 10394
rect 17119 10374 17122 10380
rect 17148 10374 17151 10400
rect 20017 10374 20020 10400
rect 20046 10394 20049 10400
rect 20693 10394 20707 10448
rect 23008 10446 23014 10448
rect 23031 10446 23037 10463
rect 23008 10443 23037 10446
rect 23099 10442 23102 10468
rect 23128 10442 23131 10468
rect 23330 10463 23359 10466
rect 23330 10446 23336 10463
rect 23353 10446 23359 10463
rect 23330 10443 23359 10446
rect 23376 10463 23405 10466
rect 23376 10446 23382 10463
rect 23399 10462 23405 10463
rect 23513 10462 23516 10468
rect 23399 10448 23516 10462
rect 23399 10446 23405 10448
rect 23376 10443 23405 10446
rect 23338 10428 23352 10443
rect 23513 10442 23516 10448
rect 23542 10442 23545 10468
rect 23974 10463 24003 10466
rect 23974 10446 23980 10463
rect 23997 10446 24003 10463
rect 23974 10443 24003 10446
rect 24020 10463 24049 10466
rect 24020 10446 24026 10463
rect 24043 10462 24049 10463
rect 24779 10463 24808 10466
rect 24779 10462 24785 10463
rect 24043 10448 24785 10462
rect 24043 10446 24049 10448
rect 24020 10443 24049 10446
rect 24779 10446 24785 10448
rect 24802 10462 24808 10463
rect 24893 10462 24896 10468
rect 24802 10448 24896 10462
rect 24802 10446 24808 10448
rect 24779 10443 24808 10446
rect 23982 10428 23996 10443
rect 24893 10442 24896 10448
rect 24922 10442 24925 10468
rect 25523 10462 25537 10550
rect 27607 10544 27610 10570
rect 27636 10564 27639 10570
rect 28389 10564 28392 10570
rect 27636 10550 28392 10564
rect 27636 10544 27639 10550
rect 28389 10544 28392 10550
rect 28418 10544 28421 10570
rect 26687 10530 26690 10536
rect 26115 10516 26690 10530
rect 25653 10497 25682 10500
rect 25653 10480 25659 10497
rect 25676 10496 25682 10497
rect 25676 10482 25974 10496
rect 25676 10480 25682 10482
rect 25653 10477 25682 10480
rect 25960 10466 25974 10482
rect 26115 10472 26129 10516
rect 26687 10510 26690 10516
rect 26716 10510 26719 10536
rect 26273 10496 26276 10502
rect 26175 10482 26276 10496
rect 26105 10469 26134 10472
rect 25906 10463 25935 10466
rect 25906 10462 25912 10463
rect 25523 10448 25912 10462
rect 25906 10446 25912 10448
rect 25929 10446 25935 10463
rect 25960 10463 25992 10466
rect 25960 10448 25969 10463
rect 25906 10443 25935 10446
rect 25963 10446 25969 10448
rect 25986 10446 25992 10463
rect 25963 10443 25992 10446
rect 26043 10442 26046 10468
rect 26072 10466 26075 10468
rect 26072 10463 26086 10466
rect 26080 10446 26086 10463
rect 26105 10452 26111 10469
rect 26128 10452 26134 10469
rect 26175 10464 26189 10482
rect 26273 10476 26276 10482
rect 26302 10476 26305 10502
rect 26871 10496 26874 10502
rect 26420 10482 26874 10496
rect 26227 10466 26230 10468
rect 26105 10449 26134 10452
rect 26167 10461 26196 10464
rect 26072 10443 26086 10446
rect 26167 10444 26173 10461
rect 26190 10444 26196 10461
rect 26072 10442 26075 10443
rect 26167 10441 26196 10444
rect 26218 10463 26230 10466
rect 26218 10446 26224 10463
rect 26256 10462 26259 10468
rect 26420 10462 26434 10482
rect 26871 10476 26874 10482
rect 26900 10496 26903 10502
rect 26900 10482 27584 10496
rect 26900 10476 26903 10482
rect 26256 10448 26434 10462
rect 26218 10443 26230 10446
rect 26227 10442 26230 10443
rect 26256 10442 26259 10448
rect 27515 10442 27518 10468
rect 27544 10442 27547 10468
rect 27570 10462 27584 10482
rect 28941 10476 28944 10502
rect 28970 10476 28973 10502
rect 28896 10463 28925 10466
rect 28896 10462 28902 10463
rect 27570 10448 28902 10462
rect 28896 10446 28902 10448
rect 28919 10446 28925 10463
rect 28896 10443 28925 10446
rect 28987 10442 28990 10468
rect 29016 10466 29019 10468
rect 29016 10443 29020 10466
rect 29016 10442 29019 10443
rect 24825 10429 24854 10432
rect 24825 10428 24831 10429
rect 23338 10414 23996 10428
rect 20046 10380 20707 10394
rect 23982 10394 23996 10414
rect 24672 10414 24831 10428
rect 24672 10400 24686 10414
rect 24825 10412 24831 10414
rect 24848 10412 24854 10429
rect 24825 10409 24854 10412
rect 27561 10408 27564 10434
rect 27590 10428 27593 10434
rect 27745 10432 27748 10434
rect 27676 10429 27705 10432
rect 27676 10428 27682 10429
rect 27590 10414 27682 10428
rect 27590 10408 27593 10414
rect 27676 10412 27682 10414
rect 27699 10412 27705 10429
rect 27676 10409 27705 10412
rect 27727 10429 27748 10432
rect 27727 10412 27733 10429
rect 27727 10409 27748 10412
rect 27745 10408 27748 10409
rect 27774 10408 27777 10434
rect 28551 10429 28580 10432
rect 28551 10412 28557 10429
rect 28574 10428 28580 10429
rect 28804 10429 28833 10432
rect 28804 10428 28810 10429
rect 28574 10414 28810 10428
rect 28574 10412 28580 10414
rect 28551 10409 28580 10412
rect 28804 10412 28810 10414
rect 28827 10412 28833 10429
rect 28804 10409 28833 10412
rect 28942 10429 28971 10432
rect 28942 10412 28948 10429
rect 28965 10428 28971 10429
rect 29125 10428 29128 10434
rect 28965 10414 29128 10428
rect 28965 10412 28971 10414
rect 28942 10409 28971 10412
rect 29125 10408 29128 10414
rect 29154 10408 29157 10434
rect 24157 10394 24160 10400
rect 23982 10380 24160 10394
rect 20046 10374 20049 10380
rect 24157 10374 24160 10380
rect 24186 10374 24189 10400
rect 24663 10374 24666 10400
rect 24692 10374 24695 10400
rect 26136 10395 26165 10398
rect 26136 10378 26142 10395
rect 26159 10394 26165 10395
rect 27147 10394 27150 10400
rect 26159 10380 27150 10394
rect 26159 10378 26165 10380
rect 26136 10375 26165 10378
rect 27147 10374 27150 10380
rect 27176 10374 27179 10400
rect 3036 10312 29992 10360
rect 7597 10272 7600 10298
rect 7626 10292 7629 10298
rect 8149 10292 8152 10298
rect 7626 10278 8152 10292
rect 7626 10272 7629 10278
rect 8149 10272 8152 10278
rect 8178 10292 8181 10298
rect 9575 10292 9578 10298
rect 8178 10278 9578 10292
rect 8178 10272 8181 10278
rect 9575 10272 9578 10278
rect 9604 10272 9607 10298
rect 14313 10272 14316 10298
rect 14342 10292 14345 10298
rect 14342 10278 15946 10292
rect 14342 10272 14345 10278
rect 9023 10238 9026 10264
rect 9052 10238 9055 10264
rect 9584 10258 9598 10272
rect 10541 10258 10544 10264
rect 9584 10244 9913 10258
rect 10281 10244 10544 10258
rect 10541 10238 10544 10244
rect 10570 10238 10573 10264
rect 14448 10259 14477 10262
rect 14448 10242 14454 10259
rect 14471 10258 14477 10259
rect 14773 10258 14776 10264
rect 14471 10244 14776 10258
rect 14471 10242 14477 10244
rect 14448 10239 14477 10242
rect 14773 10238 14776 10244
rect 14802 10238 14805 10264
rect 15740 10259 15769 10262
rect 15740 10242 15746 10259
rect 15763 10258 15769 10259
rect 15877 10258 15880 10264
rect 15763 10244 15880 10258
rect 15763 10242 15769 10244
rect 15740 10239 15769 10242
rect 15877 10238 15880 10244
rect 15906 10238 15909 10264
rect 15932 10258 15946 10278
rect 22823 10272 22826 10298
rect 22852 10292 22855 10298
rect 24111 10292 24114 10298
rect 22852 10278 24114 10292
rect 22852 10272 22855 10278
rect 24111 10272 24114 10278
rect 24140 10272 24143 10298
rect 26043 10272 26046 10298
rect 26072 10292 26075 10298
rect 26389 10293 26418 10296
rect 26389 10292 26395 10293
rect 26072 10278 26395 10292
rect 26072 10272 26075 10278
rect 26389 10276 26395 10278
rect 26412 10276 26418 10293
rect 26389 10273 26418 10276
rect 29125 10272 29128 10298
rect 29154 10296 29157 10298
rect 29154 10293 29178 10296
rect 29154 10276 29155 10293
rect 29172 10276 29178 10293
rect 29154 10273 29178 10276
rect 29154 10272 29157 10273
rect 15932 10244 15985 10258
rect 16245 10238 16248 10264
rect 16274 10238 16277 10264
rect 25583 10262 25586 10264
rect 25565 10259 25586 10262
rect 25565 10242 25571 10259
rect 25565 10239 25586 10242
rect 25583 10238 25586 10239
rect 25612 10238 25615 10264
rect 28343 10262 28346 10264
rect 28325 10259 28346 10262
rect 28325 10242 28331 10259
rect 28325 10239 28346 10242
rect 28343 10238 28346 10239
rect 28372 10238 28375 10264
rect 8058 10225 8087 10228
rect 8058 10208 8064 10225
rect 8081 10224 8087 10225
rect 8379 10224 8382 10230
rect 8081 10210 8382 10224
rect 8081 10208 8087 10210
rect 8058 10205 8087 10208
rect 8379 10204 8382 10210
rect 8408 10204 8411 10230
rect 8839 10204 8842 10230
rect 8868 10204 8871 10230
rect 8931 10204 8934 10230
rect 8960 10204 8963 10230
rect 9529 10204 9532 10230
rect 9558 10204 9561 10230
rect 15602 10225 15631 10228
rect 15602 10224 15608 10225
rect 14322 10210 15608 10224
rect 7505 10170 7508 10196
rect 7534 10190 7537 10196
rect 8012 10191 8041 10194
rect 8012 10190 8018 10191
rect 7534 10176 8018 10190
rect 7534 10170 7537 10176
rect 8012 10174 8018 10176
rect 8035 10174 8041 10191
rect 8012 10171 8041 10174
rect 9667 10170 9670 10196
rect 9696 10170 9699 10196
rect 9713 10170 9716 10196
rect 9742 10190 9745 10196
rect 10542 10191 10571 10194
rect 10542 10190 10548 10191
rect 9742 10176 10548 10190
rect 9742 10170 9745 10176
rect 10542 10174 10548 10176
rect 10565 10174 10571 10191
rect 10542 10171 10571 10174
rect 14037 10170 14040 10196
rect 14066 10190 14069 10196
rect 14322 10194 14336 10210
rect 15602 10208 15608 10210
rect 15625 10208 15631 10225
rect 15602 10205 15631 10208
rect 14314 10191 14343 10194
rect 14314 10190 14320 10191
rect 14066 10176 14320 10190
rect 14066 10170 14069 10176
rect 14314 10174 14320 10176
rect 14337 10174 14343 10191
rect 15610 10190 15624 10205
rect 25353 10204 25356 10230
rect 25382 10204 25385 10230
rect 25515 10225 25544 10228
rect 25515 10208 25521 10225
rect 25538 10224 25544 10225
rect 25675 10224 25678 10230
rect 25538 10210 25678 10224
rect 25538 10208 25544 10210
rect 25515 10205 25544 10208
rect 25675 10204 25678 10210
rect 25704 10204 25707 10230
rect 27607 10204 27610 10230
rect 27636 10224 27639 10230
rect 27975 10224 27978 10230
rect 27636 10210 27978 10224
rect 27636 10204 27639 10210
rect 27975 10204 27978 10210
rect 28004 10224 28007 10230
rect 28113 10224 28116 10230
rect 28004 10210 28116 10224
rect 28004 10204 28007 10210
rect 28113 10204 28116 10210
rect 28142 10204 28145 10230
rect 28275 10225 28304 10228
rect 28275 10208 28281 10225
rect 28298 10224 28304 10225
rect 28389 10224 28392 10230
rect 28298 10210 28392 10224
rect 28298 10208 28304 10210
rect 28275 10205 28304 10208
rect 28389 10204 28392 10210
rect 28418 10204 28421 10230
rect 15969 10190 15972 10196
rect 15610 10176 15972 10190
rect 14314 10171 14343 10174
rect 15969 10170 15972 10176
rect 15998 10170 16001 10196
rect 16614 10191 16643 10194
rect 16614 10174 16620 10191
rect 16637 10190 16643 10191
rect 17211 10190 17214 10196
rect 16637 10176 17214 10190
rect 16637 10174 16643 10176
rect 16614 10171 16643 10174
rect 17211 10170 17214 10176
rect 17240 10170 17243 10196
rect 7919 10102 7922 10128
rect 7948 10122 7951 10128
rect 8196 10123 8225 10126
rect 8196 10122 8202 10123
rect 7948 10108 8202 10122
rect 7948 10102 7951 10108
rect 8196 10106 8202 10108
rect 8219 10106 8225 10123
rect 8196 10103 8225 10106
rect 14635 10102 14638 10128
rect 14664 10122 14667 10128
rect 14865 10122 14868 10128
rect 14664 10108 14868 10122
rect 14664 10102 14667 10108
rect 14865 10102 14868 10108
rect 14894 10122 14897 10128
rect 15004 10123 15033 10126
rect 15004 10122 15010 10123
rect 14894 10108 15010 10122
rect 14894 10102 14897 10108
rect 15004 10106 15010 10108
rect 15027 10106 15033 10123
rect 15004 10103 15033 10106
rect 3036 10040 29992 10088
rect 7505 10000 7508 10026
rect 7534 10000 7537 10026
rect 9116 10021 9145 10024
rect 9116 10004 9122 10021
rect 9139 10020 9145 10021
rect 9139 10006 9460 10020
rect 9139 10004 9145 10006
rect 9116 10001 9145 10004
rect 8894 9972 9230 9986
rect 8894 9958 8908 9972
rect 7919 9932 7922 9958
rect 7948 9932 7951 9958
rect 8425 9932 8428 9958
rect 8454 9952 8457 9958
rect 8794 9953 8823 9956
rect 8794 9952 8800 9953
rect 8454 9938 8800 9952
rect 8454 9932 8457 9938
rect 8794 9936 8800 9938
rect 8817 9952 8823 9953
rect 8885 9952 8888 9958
rect 8817 9938 8888 9952
rect 8817 9936 8823 9938
rect 8794 9933 8823 9936
rect 8885 9932 8888 9938
rect 8914 9932 8917 9958
rect 9216 9956 9230 9972
rect 9208 9953 9237 9956
rect 9208 9936 9214 9953
rect 9231 9936 9237 9953
rect 9208 9933 9237 9936
rect 7460 9919 7489 9922
rect 7460 9902 7466 9919
rect 7483 9902 7489 9919
rect 7460 9899 7489 9902
rect 7468 9884 7482 9899
rect 7551 9898 7554 9924
rect 7580 9898 7583 9924
rect 7597 9898 7600 9924
rect 7626 9918 7629 9924
rect 7782 9919 7811 9922
rect 7782 9918 7788 9919
rect 7626 9904 7788 9918
rect 7626 9898 7629 9904
rect 7782 9902 7788 9904
rect 7805 9902 7811 9919
rect 7782 9899 7811 9902
rect 8977 9898 8980 9924
rect 9006 9918 9009 9924
rect 9162 9919 9191 9922
rect 9162 9918 9168 9919
rect 9006 9904 9168 9918
rect 9006 9898 9009 9904
rect 9162 9902 9168 9904
rect 9185 9918 9191 9919
rect 9253 9918 9256 9924
rect 9185 9904 9256 9918
rect 9185 9902 9191 9904
rect 9162 9899 9191 9902
rect 9253 9898 9256 9904
rect 9282 9898 9285 9924
rect 9446 9918 9460 10006
rect 9667 10000 9670 10026
rect 9696 10000 9699 10026
rect 9529 9966 9532 9992
rect 9558 9986 9561 9992
rect 9558 9972 10196 9986
rect 9558 9966 9561 9972
rect 9575 9932 9578 9958
rect 9604 9932 9607 9958
rect 10182 9956 10196 9972
rect 15969 9966 15972 9992
rect 15998 9986 16001 9992
rect 15998 9972 18476 9986
rect 15998 9966 16001 9972
rect 10174 9953 10203 9956
rect 10174 9936 10180 9953
rect 10197 9936 10203 9953
rect 10174 9933 10203 9936
rect 14360 9953 14389 9956
rect 14360 9936 14366 9953
rect 14383 9952 14389 9953
rect 14498 9953 14527 9956
rect 14383 9938 14474 9952
rect 14383 9936 14389 9938
rect 14360 9933 14389 9936
rect 9530 9919 9559 9922
rect 9530 9918 9536 9919
rect 9446 9904 9536 9918
rect 9530 9902 9536 9904
rect 9553 9918 9559 9919
rect 9713 9918 9716 9924
rect 9553 9904 9716 9918
rect 9553 9902 9559 9904
rect 9530 9899 9559 9902
rect 9713 9898 9716 9904
rect 9742 9898 9745 9924
rect 14405 9898 14408 9924
rect 14434 9898 14437 9924
rect 14460 9918 14474 9938
rect 14498 9936 14504 9953
rect 14521 9952 14527 9953
rect 15095 9952 15098 9958
rect 14521 9938 15098 9952
rect 14521 9936 14527 9938
rect 14498 9933 14527 9936
rect 15095 9932 15098 9938
rect 15124 9932 15127 9958
rect 17488 9953 17517 9956
rect 17488 9936 17494 9953
rect 17511 9952 17517 9953
rect 17901 9952 17904 9958
rect 17511 9938 17904 9952
rect 17511 9936 17517 9938
rect 17488 9933 17517 9936
rect 17901 9932 17904 9938
rect 17930 9932 17933 9958
rect 17994 9953 18023 9956
rect 17994 9936 18000 9953
rect 18017 9952 18023 9953
rect 18315 9952 18318 9958
rect 18017 9938 18318 9952
rect 18017 9936 18023 9938
rect 17994 9933 18023 9936
rect 18315 9932 18318 9938
rect 18344 9932 18347 9958
rect 14635 9918 14638 9924
rect 14460 9904 14638 9918
rect 14635 9898 14638 9904
rect 14664 9898 14667 9924
rect 17119 9898 17122 9924
rect 17148 9898 17151 9924
rect 17211 9898 17214 9924
rect 17240 9918 17243 9924
rect 17350 9919 17379 9922
rect 17350 9918 17356 9919
rect 17240 9904 17356 9918
rect 17240 9898 17243 9904
rect 17350 9902 17356 9904
rect 17373 9902 17379 9919
rect 17350 9899 17379 9902
rect 17855 9898 17858 9924
rect 17884 9898 17887 9924
rect 18462 9922 18476 9972
rect 19051 9966 19054 9992
rect 19080 9986 19083 9992
rect 19144 9987 19173 9990
rect 19144 9986 19150 9987
rect 19080 9972 19150 9986
rect 19080 9966 19083 9972
rect 19144 9970 19150 9972
rect 19167 9986 19173 9987
rect 23099 9986 23102 9992
rect 19167 9972 23102 9986
rect 19167 9970 19173 9972
rect 19144 9967 19173 9970
rect 23099 9966 23102 9972
rect 23128 9966 23131 9992
rect 22272 9953 22301 9956
rect 22272 9936 22278 9953
rect 22295 9952 22301 9953
rect 22639 9952 22642 9958
rect 22295 9938 22642 9952
rect 22295 9936 22301 9938
rect 22272 9933 22301 9936
rect 22639 9932 22642 9938
rect 22668 9932 22671 9958
rect 18454 9919 18483 9922
rect 18454 9902 18460 9919
rect 18477 9918 18483 9919
rect 19327 9918 19330 9924
rect 18477 9904 19330 9918
rect 18477 9902 18483 9904
rect 18454 9899 18483 9902
rect 19327 9898 19330 9904
rect 19356 9898 19359 9924
rect 22502 9919 22531 9922
rect 22502 9902 22508 9919
rect 22525 9918 22531 9919
rect 22685 9918 22688 9924
rect 22525 9904 22688 9918
rect 22525 9902 22531 9904
rect 22502 9899 22531 9902
rect 22685 9898 22688 9904
rect 22714 9898 22717 9924
rect 7873 9884 7876 9890
rect 7468 9870 7876 9884
rect 7873 9864 7876 9870
rect 7902 9864 7905 9890
rect 8149 9864 8152 9890
rect 8178 9864 8181 9890
rect 9024 9885 9053 9888
rect 9024 9868 9030 9885
rect 9047 9884 9053 9885
rect 9047 9870 9184 9884
rect 9047 9868 9053 9870
rect 9024 9865 9053 9868
rect 9069 9830 9072 9856
rect 9098 9830 9101 9856
rect 9170 9850 9184 9870
rect 10311 9864 10314 9890
rect 10340 9864 10343 9890
rect 10541 9864 10544 9890
rect 10570 9864 10573 9890
rect 10817 9864 10820 9890
rect 10846 9864 10849 9890
rect 13899 9884 13902 9890
rect 10925 9870 13902 9884
rect 13899 9864 13902 9870
rect 13928 9864 13931 9890
rect 14498 9885 14527 9888
rect 14498 9868 14504 9885
rect 14521 9884 14527 9885
rect 14589 9884 14592 9890
rect 14521 9870 14592 9884
rect 14521 9868 14527 9870
rect 14498 9865 14527 9868
rect 14589 9864 14592 9870
rect 14618 9864 14621 9890
rect 18577 9885 18606 9888
rect 18577 9884 18583 9885
rect 18278 9870 18583 9884
rect 9989 9850 9992 9856
rect 9170 9836 9992 9850
rect 9989 9830 9992 9836
rect 10018 9850 10021 9856
rect 11048 9851 11077 9854
rect 11048 9850 11054 9851
rect 10018 9836 11054 9850
rect 10018 9830 10021 9836
rect 11048 9834 11054 9836
rect 11071 9834 11077 9851
rect 11048 9831 11077 9834
rect 15233 9830 15236 9856
rect 15262 9850 15265 9856
rect 17166 9851 17195 9854
rect 17166 9850 17172 9851
rect 15262 9836 17172 9850
rect 15262 9830 15265 9836
rect 17166 9834 17172 9836
rect 17189 9834 17195 9851
rect 17166 9831 17195 9834
rect 17856 9851 17885 9854
rect 17856 9834 17862 9851
rect 17879 9850 17885 9851
rect 18278 9850 18292 9870
rect 18577 9868 18583 9870
rect 18600 9868 18606 9885
rect 18577 9865 18606 9868
rect 22317 9864 22320 9890
rect 22346 9864 22349 9890
rect 22547 9864 22550 9890
rect 22576 9864 22579 9890
rect 22594 9885 22623 9888
rect 22594 9868 22600 9885
rect 22617 9884 22623 9885
rect 22731 9884 22734 9890
rect 22617 9870 22734 9884
rect 22617 9868 22623 9870
rect 22594 9865 22623 9868
rect 22731 9864 22734 9870
rect 22760 9864 22763 9890
rect 17879 9836 18292 9850
rect 17879 9834 17885 9836
rect 17856 9831 17885 9834
rect 22179 9830 22182 9856
rect 22208 9850 22211 9856
rect 22326 9850 22340 9864
rect 27239 9850 27242 9856
rect 22208 9836 27242 9850
rect 22208 9830 22211 9836
rect 27239 9830 27242 9836
rect 27268 9830 27271 9856
rect 28481 9830 28484 9856
rect 28510 9850 28513 9856
rect 28619 9850 28622 9856
rect 28510 9836 28622 9850
rect 28510 9830 28513 9836
rect 28619 9830 28622 9836
rect 28648 9830 28651 9856
rect 3036 9768 29992 9816
rect 8885 9728 8888 9754
rect 8914 9728 8917 9754
rect 8978 9749 9007 9752
rect 8978 9732 8984 9749
rect 9001 9732 9007 9749
rect 8978 9729 9007 9732
rect 7873 9694 7876 9720
rect 7902 9714 7905 9720
rect 8103 9714 8106 9720
rect 7902 9700 8106 9714
rect 7902 9694 7905 9700
rect 8103 9694 8106 9700
rect 8132 9714 8135 9720
rect 8333 9714 8336 9720
rect 8132 9700 8336 9714
rect 8132 9694 8135 9700
rect 8333 9694 8336 9700
rect 8362 9694 8365 9720
rect 8840 9715 8869 9718
rect 8840 9698 8846 9715
rect 8863 9714 8869 9715
rect 8931 9714 8934 9720
rect 8863 9700 8934 9714
rect 8863 9698 8869 9700
rect 8840 9695 8869 9698
rect 8931 9694 8934 9700
rect 8960 9694 8963 9720
rect 7551 9660 7554 9686
rect 7580 9680 7583 9686
rect 7920 9681 7949 9684
rect 7920 9680 7926 9681
rect 7580 9666 7926 9680
rect 7580 9660 7583 9666
rect 7920 9664 7926 9666
rect 7943 9680 7949 9681
rect 8342 9680 8356 9694
rect 8794 9681 8823 9684
rect 8794 9680 8800 9681
rect 7943 9666 8287 9680
rect 8342 9666 8800 9680
rect 7943 9664 7949 9666
rect 7920 9661 7949 9664
rect 7873 9626 7876 9652
rect 7902 9626 7905 9652
rect 8273 9646 8287 9666
rect 8794 9664 8800 9666
rect 8817 9664 8823 9681
rect 8986 9680 9000 9729
rect 14405 9728 14408 9754
rect 14434 9748 14437 9754
rect 14452 9749 14481 9752
rect 14452 9748 14458 9749
rect 14434 9734 14458 9748
rect 14434 9728 14437 9734
rect 14452 9732 14458 9734
rect 14475 9732 14481 9749
rect 14452 9729 14481 9732
rect 20615 9728 20618 9754
rect 20644 9728 20647 9754
rect 23421 9728 23424 9754
rect 23450 9728 23453 9754
rect 9484 9715 9513 9718
rect 9484 9698 9490 9715
rect 9507 9714 9513 9715
rect 9713 9714 9716 9720
rect 9507 9700 9716 9714
rect 9507 9698 9513 9700
rect 9484 9695 9513 9698
rect 9713 9694 9716 9700
rect 9742 9694 9745 9720
rect 14360 9715 14389 9718
rect 14360 9698 14366 9715
rect 14383 9714 14389 9715
rect 15049 9714 15052 9720
rect 14383 9700 15052 9714
rect 14383 9698 14389 9700
rect 14360 9695 14389 9698
rect 15049 9694 15052 9700
rect 15078 9694 15081 9720
rect 17027 9694 17030 9720
rect 17056 9714 17059 9720
rect 17166 9715 17195 9718
rect 17166 9714 17172 9715
rect 17056 9700 17172 9714
rect 17056 9694 17059 9700
rect 17166 9698 17172 9700
rect 17189 9714 17195 9715
rect 17211 9714 17214 9720
rect 17189 9700 17214 9714
rect 17189 9698 17195 9700
rect 17166 9695 17195 9698
rect 17211 9694 17214 9700
rect 17240 9694 17243 9720
rect 19190 9715 19219 9718
rect 19190 9698 19196 9715
rect 19213 9714 19219 9715
rect 19235 9714 19238 9720
rect 19213 9700 19238 9714
rect 19213 9698 19219 9700
rect 19190 9695 19219 9698
rect 19235 9694 19238 9700
rect 19264 9694 19267 9720
rect 22317 9714 22320 9720
rect 20532 9700 22320 9714
rect 9575 9680 9578 9686
rect 8986 9666 9578 9680
rect 8794 9661 8823 9664
rect 9575 9660 9578 9666
rect 9604 9660 9607 9686
rect 9989 9660 9992 9686
rect 10018 9660 10021 9686
rect 14497 9660 14500 9686
rect 14526 9660 14529 9686
rect 17074 9681 17103 9684
rect 17074 9664 17080 9681
rect 17097 9680 17103 9681
rect 17119 9680 17122 9686
rect 17097 9666 17122 9680
rect 17097 9664 17103 9666
rect 17074 9661 17103 9664
rect 17119 9660 17122 9666
rect 17148 9660 17151 9686
rect 19097 9660 19100 9686
rect 19126 9660 19129 9686
rect 19143 9660 19146 9686
rect 19172 9660 19175 9686
rect 20532 9684 20546 9700
rect 22317 9694 22320 9700
rect 22346 9694 22349 9720
rect 22639 9694 22642 9720
rect 22668 9714 22671 9720
rect 22668 9700 23352 9714
rect 22668 9694 22671 9700
rect 20524 9681 20553 9684
rect 20524 9664 20530 9681
rect 20547 9664 20553 9681
rect 20524 9661 20553 9664
rect 20569 9660 20572 9686
rect 20598 9660 20601 9686
rect 22547 9660 22550 9686
rect 22576 9680 22579 9686
rect 22594 9681 22623 9684
rect 22594 9680 22600 9681
rect 22576 9666 22600 9680
rect 22576 9660 22579 9666
rect 22594 9664 22600 9666
rect 22617 9664 22623 9681
rect 22594 9661 22623 9664
rect 22685 9660 22688 9686
rect 22714 9660 22717 9686
rect 22731 9660 22734 9686
rect 22760 9680 22763 9686
rect 23338 9684 23352 9700
rect 25353 9694 25356 9720
rect 25382 9714 25385 9720
rect 25382 9700 25537 9714
rect 25382 9694 25385 9700
rect 23100 9681 23129 9684
rect 23100 9680 23106 9681
rect 22760 9666 23106 9680
rect 22760 9660 22763 9666
rect 23100 9664 23106 9666
rect 23123 9664 23129 9681
rect 23100 9661 23129 9664
rect 23330 9681 23359 9684
rect 23330 9664 23336 9681
rect 23353 9664 23359 9681
rect 25523 9680 25537 9700
rect 27239 9694 27242 9720
rect 27268 9714 27271 9720
rect 28987 9714 28990 9720
rect 27268 9700 28990 9714
rect 27268 9694 27271 9700
rect 28987 9694 28990 9700
rect 29016 9694 29019 9720
rect 25629 9680 25632 9686
rect 25523 9666 25632 9680
rect 23330 9661 23359 9664
rect 25629 9660 25632 9666
rect 25658 9660 25661 9686
rect 28260 9666 28504 9680
rect 8471 9646 8474 9652
rect 8273 9632 8474 9646
rect 8471 9626 8474 9632
rect 8500 9646 8503 9652
rect 8885 9646 8888 9652
rect 8500 9632 8888 9646
rect 8500 9626 8503 9632
rect 8885 9626 8888 9632
rect 8914 9646 8917 9652
rect 8978 9647 9007 9650
rect 8978 9646 8984 9647
rect 8914 9632 8984 9646
rect 8914 9626 8917 9632
rect 8978 9630 8984 9632
rect 9001 9630 9007 9647
rect 8978 9627 9007 9630
rect 9668 9647 9697 9650
rect 9668 9630 9674 9647
rect 9691 9646 9697 9647
rect 9944 9647 9973 9650
rect 9944 9646 9950 9647
rect 9691 9632 9950 9646
rect 9691 9630 9697 9632
rect 9668 9627 9697 9630
rect 9944 9630 9950 9632
rect 9967 9630 9973 9647
rect 9944 9627 9973 9630
rect 10174 9647 10203 9650
rect 10174 9630 10180 9647
rect 10197 9646 10203 9647
rect 10311 9646 10314 9652
rect 10197 9632 10314 9646
rect 10197 9630 10203 9632
rect 10174 9627 10203 9630
rect 10311 9626 10314 9632
rect 10340 9626 10343 9652
rect 16567 9626 16570 9652
rect 16596 9646 16599 9652
rect 16935 9646 16938 9652
rect 16596 9632 16938 9646
rect 16596 9626 16599 9632
rect 16935 9626 16938 9632
rect 16964 9646 16967 9652
rect 17258 9647 17287 9650
rect 17258 9646 17264 9647
rect 16964 9632 17264 9646
rect 16964 9626 16967 9632
rect 17258 9630 17264 9632
rect 17281 9630 17287 9647
rect 17258 9627 17287 9630
rect 19005 9626 19008 9652
rect 19034 9626 19037 9652
rect 19374 9647 19403 9650
rect 19374 9630 19380 9647
rect 19397 9646 19403 9647
rect 20708 9647 20737 9650
rect 19397 9632 20684 9646
rect 19397 9630 19403 9632
rect 19374 9627 19403 9630
rect 8839 9592 8842 9618
rect 8868 9592 8871 9618
rect 19879 9592 19882 9618
rect 19908 9612 19911 9618
rect 20570 9613 20599 9616
rect 20570 9612 20576 9613
rect 19908 9598 20576 9612
rect 19908 9592 19911 9598
rect 20570 9596 20576 9598
rect 20593 9596 20599 9613
rect 20670 9612 20684 9632
rect 20708 9630 20714 9647
rect 20731 9646 20737 9647
rect 22087 9646 22090 9652
rect 20731 9632 22090 9646
rect 20731 9630 20737 9632
rect 20708 9627 20737 9630
rect 22087 9626 22090 9632
rect 22116 9626 22119 9652
rect 25353 9626 25356 9652
rect 25382 9646 25385 9652
rect 28260 9646 28274 9666
rect 25382 9632 28274 9646
rect 25382 9626 25385 9632
rect 28297 9626 28300 9652
rect 28326 9646 28329 9652
rect 28435 9646 28438 9652
rect 28326 9632 28438 9646
rect 28326 9626 28329 9632
rect 28435 9626 28438 9632
rect 28464 9626 28467 9652
rect 28490 9646 28504 9666
rect 29401 9646 29404 9652
rect 28490 9632 29404 9646
rect 29401 9626 29404 9632
rect 29430 9626 29433 9652
rect 21719 9612 21722 9618
rect 20670 9598 21722 9612
rect 20570 9593 20599 9596
rect 21719 9592 21722 9598
rect 21748 9612 21751 9618
rect 24617 9612 24620 9618
rect 21748 9598 24620 9612
rect 21748 9592 21751 9598
rect 24617 9592 24620 9598
rect 24646 9592 24649 9618
rect 26963 9592 26966 9618
rect 26992 9612 26995 9618
rect 28849 9612 28852 9618
rect 26992 9598 28852 9612
rect 26992 9592 26995 9598
rect 28849 9592 28852 9598
rect 28878 9592 28881 9618
rect 7781 9558 7784 9584
rect 7810 9578 7813 9584
rect 8104 9579 8133 9582
rect 8104 9578 8110 9579
rect 7810 9564 8110 9578
rect 7810 9558 7813 9564
rect 8104 9562 8110 9564
rect 8127 9562 8133 9579
rect 8104 9559 8133 9562
rect 14359 9558 14362 9584
rect 14388 9558 14391 9584
rect 25859 9558 25862 9584
rect 25888 9578 25891 9584
rect 28665 9578 28668 9584
rect 25888 9564 28668 9578
rect 25888 9558 25891 9564
rect 28665 9558 28668 9564
rect 28694 9558 28697 9584
rect 3036 9496 29992 9544
rect 15049 9456 15052 9482
rect 15078 9456 15081 9482
rect 20524 9477 20553 9480
rect 20524 9460 20530 9477
rect 20547 9476 20553 9477
rect 20569 9476 20572 9482
rect 20547 9462 20572 9476
rect 20547 9460 20553 9462
rect 20524 9457 20553 9460
rect 20569 9456 20572 9462
rect 20598 9456 20601 9482
rect 23973 9456 23976 9482
rect 24002 9476 24005 9482
rect 26687 9476 26690 9482
rect 24002 9462 26690 9476
rect 24002 9456 24005 9462
rect 26687 9456 26690 9462
rect 26716 9456 26719 9482
rect 26733 9456 26736 9482
rect 26762 9476 26765 9482
rect 27010 9477 27039 9480
rect 27010 9476 27016 9477
rect 26762 9462 27016 9476
rect 26762 9456 26765 9462
rect 27010 9460 27016 9462
rect 27033 9460 27039 9477
rect 29033 9476 29036 9482
rect 27010 9457 27039 9460
rect 28973 9462 29036 9476
rect 21397 9422 21400 9448
rect 21426 9442 21429 9448
rect 23881 9442 23884 9448
rect 21426 9428 23884 9442
rect 21426 9422 21429 9428
rect 23881 9422 23884 9428
rect 23910 9422 23913 9448
rect 7781 9388 7784 9414
rect 7810 9388 7813 9414
rect 8656 9409 8685 9412
rect 8656 9392 8662 9409
rect 8679 9408 8685 9409
rect 8885 9408 8888 9414
rect 8679 9394 8888 9408
rect 8679 9392 8685 9394
rect 8656 9389 8685 9392
rect 8885 9388 8888 9394
rect 8914 9388 8917 9414
rect 15004 9409 15033 9412
rect 15004 9408 15010 9409
rect 14552 9394 15010 9408
rect 7597 9354 7600 9380
rect 7626 9374 7629 9380
rect 7644 9375 7673 9378
rect 7644 9374 7650 9375
rect 7626 9360 7650 9374
rect 7626 9354 7629 9360
rect 7644 9358 7650 9360
rect 7667 9358 7673 9375
rect 7644 9355 7673 9358
rect 14037 9354 14040 9380
rect 14066 9354 14069 9380
rect 14172 9375 14201 9378
rect 14172 9358 14178 9375
rect 14195 9374 14201 9375
rect 14359 9374 14362 9380
rect 14195 9360 14362 9374
rect 14195 9358 14201 9360
rect 14172 9355 14201 9358
rect 14359 9354 14362 9360
rect 14388 9354 14391 9380
rect 14405 9354 14408 9380
rect 14434 9374 14437 9380
rect 14552 9374 14566 9394
rect 15004 9392 15010 9394
rect 15027 9392 15033 9409
rect 15004 9389 15033 9392
rect 15095 9388 15098 9414
rect 15124 9388 15127 9414
rect 19005 9388 19008 9414
rect 19034 9408 19037 9414
rect 21351 9408 21354 9414
rect 19034 9394 19626 9408
rect 19034 9388 19037 9394
rect 19612 9380 19626 9394
rect 20624 9394 21354 9408
rect 14958 9375 14987 9378
rect 14958 9374 14964 9375
rect 14434 9360 14566 9374
rect 14736 9360 14964 9374
rect 14434 9354 14437 9360
rect 7735 9320 7738 9346
rect 7764 9340 7767 9346
rect 7764 9326 8027 9340
rect 7764 9320 7767 9326
rect 8149 9320 8152 9346
rect 8178 9320 8181 9346
rect 14543 9286 14546 9312
rect 14572 9306 14575 9312
rect 14736 9310 14750 9360
rect 14958 9358 14964 9360
rect 14981 9358 14987 9375
rect 14958 9355 14987 9358
rect 15878 9375 15907 9378
rect 15878 9358 15884 9375
rect 15901 9374 15907 9375
rect 16107 9374 16110 9380
rect 15901 9360 16110 9374
rect 15901 9358 15907 9360
rect 15878 9355 15907 9358
rect 16107 9354 16110 9360
rect 16136 9354 16139 9380
rect 18637 9354 18640 9380
rect 18666 9374 18669 9380
rect 18868 9375 18897 9378
rect 18868 9374 18874 9375
rect 18666 9360 18874 9374
rect 18666 9354 18669 9360
rect 18868 9358 18874 9360
rect 18891 9358 18897 9375
rect 18868 9355 18897 9358
rect 18960 9375 18989 9378
rect 18960 9358 18966 9375
rect 18983 9374 18989 9375
rect 19097 9374 19100 9380
rect 18983 9360 19100 9374
rect 18983 9358 18989 9360
rect 18960 9355 18989 9358
rect 19097 9354 19100 9360
rect 19126 9374 19129 9380
rect 19281 9374 19284 9380
rect 19126 9360 19284 9374
rect 19126 9354 19129 9360
rect 19281 9354 19284 9360
rect 19310 9354 19313 9380
rect 19374 9375 19403 9378
rect 19374 9358 19380 9375
rect 19397 9358 19403 9375
rect 19374 9355 19403 9358
rect 15463 9320 15466 9346
rect 15492 9340 15495 9346
rect 15740 9341 15769 9344
rect 15740 9340 15746 9341
rect 15492 9326 15746 9340
rect 15492 9320 15495 9326
rect 15740 9324 15746 9326
rect 15763 9324 15769 9341
rect 15740 9321 15769 9324
rect 15832 9341 15861 9344
rect 15832 9324 15838 9341
rect 15855 9340 15861 9341
rect 15855 9326 15900 9340
rect 15855 9324 15861 9326
rect 15832 9321 15861 9324
rect 15886 9312 15900 9326
rect 19143 9320 19146 9346
rect 19172 9340 19175 9346
rect 19382 9340 19396 9355
rect 19603 9354 19606 9380
rect 19632 9354 19635 9380
rect 20247 9354 20250 9380
rect 20276 9374 20279 9380
rect 20624 9378 20638 9394
rect 21351 9388 21354 9394
rect 21380 9388 21383 9414
rect 22179 9408 22182 9414
rect 22096 9394 22182 9408
rect 20616 9375 20645 9378
rect 20616 9374 20622 9375
rect 20276 9360 20622 9374
rect 20276 9354 20279 9360
rect 20616 9358 20622 9360
rect 20639 9358 20645 9375
rect 20616 9355 20645 9358
rect 20661 9354 20664 9380
rect 20690 9354 20693 9380
rect 20726 9375 20755 9378
rect 20726 9358 20732 9375
rect 20749 9374 20755 9375
rect 22096 9374 22110 9394
rect 22179 9388 22182 9394
rect 22208 9388 22211 9414
rect 22547 9408 22550 9414
rect 22234 9394 22550 9408
rect 22234 9378 22248 9394
rect 22547 9388 22550 9394
rect 22576 9408 22579 9414
rect 22777 9408 22780 9414
rect 22576 9394 22780 9408
rect 22576 9388 22579 9394
rect 22777 9388 22780 9394
rect 22806 9388 22809 9414
rect 23237 9388 23240 9414
rect 23266 9408 23269 9414
rect 23835 9408 23838 9414
rect 23266 9394 23838 9408
rect 23266 9388 23269 9394
rect 23835 9388 23838 9394
rect 23864 9408 23867 9414
rect 23974 9409 24003 9412
rect 23974 9408 23980 9409
rect 23864 9394 23980 9408
rect 23864 9388 23867 9394
rect 23974 9392 23980 9394
rect 23997 9392 24003 9409
rect 23974 9389 24003 9392
rect 25261 9388 25264 9414
rect 25290 9388 25293 9414
rect 27055 9408 27058 9414
rect 26880 9394 27058 9408
rect 26880 9380 26894 9394
rect 27055 9388 27058 9394
rect 27084 9388 27087 9414
rect 27147 9388 27150 9414
rect 27176 9388 27179 9414
rect 27975 9388 27978 9414
rect 28004 9388 28007 9414
rect 20749 9360 22110 9374
rect 22134 9375 22163 9378
rect 20749 9358 20755 9360
rect 20726 9355 20755 9358
rect 22134 9358 22140 9375
rect 22157 9358 22163 9375
rect 22134 9355 22163 9358
rect 22226 9375 22255 9378
rect 22226 9358 22232 9375
rect 22249 9358 22255 9375
rect 22226 9355 22255 9358
rect 20431 9340 20434 9346
rect 19172 9326 20434 9340
rect 19172 9320 19175 9326
rect 20431 9320 20434 9326
rect 20460 9320 20463 9346
rect 20523 9320 20526 9346
rect 20552 9320 20555 9346
rect 21995 9320 21998 9346
rect 22024 9340 22027 9346
rect 22142 9340 22156 9355
rect 22639 9354 22642 9380
rect 22668 9354 22671 9380
rect 22685 9354 22688 9380
rect 22714 9374 22717 9380
rect 22870 9375 22899 9378
rect 22870 9374 22876 9375
rect 22714 9360 22876 9374
rect 22714 9354 22717 9360
rect 22870 9358 22876 9360
rect 22893 9358 22899 9375
rect 22870 9355 22899 9358
rect 23421 9354 23424 9380
rect 23450 9374 23453 9380
rect 25449 9375 25478 9378
rect 25449 9374 25455 9375
rect 23450 9360 25455 9374
rect 23450 9354 23453 9360
rect 25449 9358 25455 9360
rect 25472 9374 25478 9375
rect 26871 9374 26874 9380
rect 25472 9360 26874 9374
rect 25472 9358 25478 9360
rect 25449 9355 25478 9358
rect 26871 9354 26874 9360
rect 26900 9354 26903 9380
rect 26964 9375 26993 9378
rect 26964 9358 26970 9375
rect 26987 9374 26993 9375
rect 28973 9374 28987 9462
rect 29033 9456 29036 9462
rect 29062 9456 29065 9482
rect 29493 9456 29496 9482
rect 29522 9456 29525 9482
rect 26987 9360 28987 9374
rect 26987 9358 26993 9360
rect 26964 9355 26993 9358
rect 29171 9354 29174 9380
rect 29200 9374 29203 9380
rect 29585 9374 29588 9380
rect 29200 9360 29588 9374
rect 29200 9354 29203 9360
rect 29585 9354 29588 9360
rect 29614 9354 29617 9380
rect 29677 9354 29680 9380
rect 29706 9378 29709 9380
rect 29706 9374 29710 9378
rect 29706 9360 29728 9374
rect 29706 9355 29710 9360
rect 29706 9354 29709 9355
rect 24203 9344 24206 9346
rect 24134 9341 24163 9344
rect 24134 9340 24140 9341
rect 22024 9326 22156 9340
rect 24028 9326 24140 9340
rect 22024 9320 22027 9326
rect 14728 9307 14757 9310
rect 14728 9306 14734 9307
rect 14572 9292 14734 9306
rect 14572 9286 14575 9292
rect 14728 9290 14734 9292
rect 14751 9290 14757 9307
rect 14728 9287 14757 9290
rect 15785 9286 15788 9312
rect 15814 9286 15817 9312
rect 15877 9286 15880 9312
rect 15906 9286 15909 9312
rect 18959 9286 18962 9312
rect 18988 9306 18991 9312
rect 19052 9307 19081 9310
rect 19052 9306 19058 9307
rect 18988 9292 19058 9306
rect 18988 9286 18991 9292
rect 19052 9290 19058 9292
rect 19075 9290 19081 9307
rect 19052 9287 19081 9290
rect 19696 9307 19725 9310
rect 19696 9290 19702 9307
rect 19719 9306 19725 9307
rect 21949 9306 21952 9312
rect 19719 9292 21952 9306
rect 19719 9290 19725 9292
rect 19696 9287 19725 9290
rect 21949 9286 21952 9292
rect 21978 9286 21981 9312
rect 22961 9286 22964 9312
rect 22990 9286 22993 9312
rect 23973 9286 23976 9312
rect 24002 9306 24005 9312
rect 24028 9306 24042 9326
rect 24134 9324 24140 9326
rect 24157 9324 24163 9341
rect 24134 9321 24163 9324
rect 24185 9341 24206 9344
rect 24185 9324 24191 9341
rect 24185 9321 24206 9324
rect 24203 9320 24206 9321
rect 24232 9320 24235 9346
rect 25009 9341 25038 9344
rect 25009 9324 25015 9341
rect 25032 9340 25038 9341
rect 25262 9341 25291 9344
rect 25262 9340 25268 9341
rect 25032 9326 25268 9340
rect 25032 9324 25038 9326
rect 25009 9321 25038 9324
rect 25262 9324 25268 9326
rect 25285 9324 25291 9341
rect 25262 9321 25291 9324
rect 25353 9320 25356 9346
rect 25382 9320 25385 9346
rect 25399 9320 25402 9346
rect 25428 9320 25431 9346
rect 28021 9320 28024 9346
rect 28050 9340 28053 9346
rect 28205 9344 28208 9346
rect 28136 9341 28165 9344
rect 28136 9340 28142 9341
rect 28050 9326 28142 9340
rect 28050 9320 28053 9326
rect 28136 9324 28142 9326
rect 28159 9324 28165 9341
rect 28136 9321 28165 9324
rect 28187 9341 28208 9344
rect 28187 9324 28193 9341
rect 28187 9321 28208 9324
rect 28205 9320 28208 9321
rect 28234 9320 28237 9346
rect 29011 9341 29040 9344
rect 29011 9324 29017 9341
rect 29034 9340 29040 9341
rect 29494 9341 29523 9344
rect 29494 9340 29500 9341
rect 29034 9326 29500 9340
rect 29034 9324 29040 9326
rect 29011 9321 29040 9324
rect 29494 9324 29500 9326
rect 29517 9324 29523 9341
rect 29494 9321 29523 9324
rect 29631 9320 29634 9346
rect 29660 9320 29663 9346
rect 24002 9292 24042 9306
rect 24002 9286 24005 9292
rect 26917 9286 26920 9312
rect 26946 9306 26949 9312
rect 27010 9307 27039 9310
rect 27010 9306 27016 9307
rect 26946 9292 27016 9306
rect 26946 9286 26949 9292
rect 27010 9290 27016 9292
rect 27033 9290 27039 9307
rect 27010 9287 27039 9290
rect 27056 9307 27085 9310
rect 27056 9290 27062 9307
rect 27079 9306 27085 9307
rect 27147 9306 27150 9312
rect 27079 9292 27150 9306
rect 27079 9290 27085 9292
rect 27056 9287 27085 9290
rect 27147 9286 27150 9292
rect 27176 9286 27179 9312
rect 3036 9224 29992 9272
rect 14497 9184 14500 9210
rect 14526 9204 14529 9210
rect 14728 9205 14757 9208
rect 14728 9204 14734 9205
rect 14526 9190 14734 9204
rect 14526 9184 14529 9190
rect 14728 9188 14734 9190
rect 14751 9188 14757 9205
rect 14728 9185 14757 9188
rect 15863 9190 17947 9204
rect 13807 9170 13810 9176
rect 13770 9156 13810 9170
rect 13770 9140 13784 9156
rect 13807 9150 13810 9156
rect 13836 9170 13839 9176
rect 14405 9170 14408 9176
rect 13836 9156 14408 9170
rect 13836 9150 13839 9156
rect 14405 9150 14408 9156
rect 14434 9150 14437 9176
rect 14635 9170 14638 9176
rect 14598 9156 14638 9170
rect 13762 9137 13791 9140
rect 13762 9120 13768 9137
rect 13785 9120 13791 9137
rect 13762 9117 13791 9120
rect 13854 9137 13883 9140
rect 13854 9120 13860 9137
rect 13877 9136 13883 9137
rect 14129 9136 14132 9142
rect 13877 9122 14132 9136
rect 13877 9120 13883 9122
rect 13854 9117 13883 9120
rect 14129 9116 14132 9122
rect 14158 9116 14161 9142
rect 14543 9116 14546 9142
rect 14572 9116 14575 9142
rect 14598 9106 14612 9156
rect 14635 9150 14638 9156
rect 14664 9170 14667 9176
rect 15863 9170 15877 9190
rect 14664 9156 15877 9170
rect 14664 9150 14667 9156
rect 15923 9150 15926 9176
rect 15952 9150 15955 9176
rect 15280 9137 15309 9140
rect 15280 9120 15286 9137
rect 15303 9136 15309 9137
rect 15932 9136 15946 9150
rect 15303 9122 15946 9136
rect 15303 9120 15309 9122
rect 15280 9117 15309 9120
rect 15969 9116 15972 9142
rect 15998 9136 16001 9142
rect 16052 9137 16081 9140
rect 16052 9136 16058 9137
rect 15998 9122 16058 9136
rect 15998 9116 16001 9122
rect 16052 9120 16058 9122
rect 16075 9120 16081 9137
rect 17933 9136 17947 9190
rect 19235 9184 19238 9210
rect 19264 9184 19267 9210
rect 20523 9184 20526 9210
rect 20552 9204 20555 9210
rect 20869 9205 20898 9208
rect 20869 9204 20875 9205
rect 20552 9190 20875 9204
rect 20552 9184 20555 9190
rect 20869 9188 20875 9190
rect 20892 9188 20898 9205
rect 20869 9185 20898 9188
rect 22593 9184 22596 9210
rect 22622 9204 22625 9210
rect 22778 9205 22807 9208
rect 22778 9204 22784 9205
rect 22622 9190 22784 9204
rect 22622 9184 22625 9190
rect 22778 9188 22784 9190
rect 22801 9188 22807 9205
rect 22778 9185 22807 9188
rect 23421 9184 23424 9210
rect 23450 9184 23453 9210
rect 24871 9205 24900 9208
rect 24871 9188 24877 9205
rect 24894 9204 24900 9205
rect 25399 9204 25402 9210
rect 24894 9190 25402 9204
rect 24894 9188 24900 9190
rect 24871 9185 24900 9188
rect 25399 9184 25402 9190
rect 25428 9184 25431 9210
rect 26917 9184 26920 9210
rect 26946 9184 26949 9210
rect 29149 9205 29178 9208
rect 29149 9188 29155 9205
rect 29172 9204 29178 9205
rect 29631 9204 29634 9210
rect 29172 9190 29634 9204
rect 29172 9188 29178 9190
rect 29149 9185 29178 9188
rect 29631 9184 29634 9190
rect 29660 9184 29663 9210
rect 18637 9150 18640 9176
rect 18666 9170 18669 9176
rect 19244 9170 19258 9184
rect 20063 9174 20066 9176
rect 19282 9171 19311 9174
rect 19282 9170 19288 9171
rect 18666 9156 19288 9170
rect 18666 9150 18669 9156
rect 19282 9154 19288 9156
rect 19305 9154 19311 9171
rect 19282 9151 19311 9154
rect 20045 9171 20066 9174
rect 20045 9154 20051 9171
rect 20092 9170 20095 9176
rect 22731 9170 22734 9176
rect 20092 9156 20178 9170
rect 20045 9151 20066 9154
rect 20063 9150 20066 9151
rect 20092 9150 20095 9156
rect 18960 9137 18989 9140
rect 18960 9136 18966 9137
rect 17933 9122 18966 9136
rect 16052 9117 16081 9120
rect 18960 9120 18966 9122
rect 18983 9136 18989 9137
rect 19143 9136 19146 9142
rect 18983 9122 19146 9136
rect 18983 9120 18989 9122
rect 18960 9117 18989 9120
rect 19143 9116 19146 9122
rect 19172 9116 19175 9142
rect 19190 9137 19219 9140
rect 19190 9120 19196 9137
rect 19213 9120 19219 9137
rect 19190 9117 19219 9120
rect 14590 9103 14619 9106
rect 14590 9102 14596 9103
rect 14552 9088 14596 9102
rect 14552 9074 14566 9088
rect 14590 9086 14596 9088
rect 14613 9086 14619 9103
rect 14590 9083 14619 9086
rect 15234 9103 15263 9106
rect 15234 9086 15240 9103
rect 15257 9086 15263 9103
rect 15234 9083 15263 9086
rect 14543 9048 14546 9074
rect 14572 9048 14575 9074
rect 14728 9069 14757 9072
rect 14728 9052 14734 9069
rect 14751 9068 14757 9069
rect 15242 9068 15256 9083
rect 15463 9082 15466 9108
rect 15492 9082 15495 9108
rect 15924 9103 15953 9106
rect 15924 9086 15930 9103
rect 15947 9086 15953 9103
rect 15924 9083 15953 9086
rect 14751 9054 15256 9068
rect 14751 9052 14757 9054
rect 14728 9049 14757 9052
rect 13762 9035 13791 9038
rect 13762 9018 13768 9035
rect 13785 9034 13791 9035
rect 14451 9034 14454 9040
rect 13785 9020 14454 9034
rect 13785 9018 13791 9020
rect 13762 9015 13791 9018
rect 14451 9014 14454 9020
rect 14480 9014 14483 9040
rect 15932 9034 15946 9083
rect 17073 9082 17076 9108
rect 17102 9082 17105 9108
rect 17119 9082 17122 9108
rect 17148 9082 17151 9108
rect 17165 9082 17168 9108
rect 17194 9102 17197 9108
rect 17212 9103 17241 9106
rect 17212 9102 17218 9103
rect 17194 9088 17218 9102
rect 17194 9082 17197 9088
rect 17212 9086 17218 9088
rect 17235 9086 17241 9103
rect 17212 9083 17241 9086
rect 18913 9082 18916 9108
rect 18942 9102 18945 9108
rect 19006 9103 19035 9106
rect 19006 9102 19012 9103
rect 18942 9088 19012 9102
rect 18942 9082 18945 9088
rect 19006 9086 19012 9088
rect 19029 9086 19035 9103
rect 19198 9102 19212 9117
rect 19235 9116 19238 9142
rect 19264 9136 19267 9142
rect 19603 9136 19606 9142
rect 19264 9122 19606 9136
rect 19264 9116 19267 9122
rect 19603 9116 19606 9122
rect 19632 9116 19635 9142
rect 19995 9137 20024 9140
rect 19995 9120 20001 9137
rect 20018 9136 20024 9137
rect 20109 9136 20112 9142
rect 20018 9122 20112 9136
rect 20018 9120 20024 9122
rect 19995 9117 20024 9120
rect 20109 9116 20112 9122
rect 20138 9116 20141 9142
rect 20164 9136 20178 9156
rect 22602 9156 22734 9170
rect 20569 9136 20572 9142
rect 20164 9122 20572 9136
rect 20569 9116 20572 9122
rect 20598 9136 20601 9142
rect 20598 9122 20707 9136
rect 20598 9116 20601 9122
rect 19198 9088 19304 9102
rect 19006 9083 19035 9086
rect 16614 9069 16643 9072
rect 16614 9052 16620 9069
rect 16637 9068 16643 9069
rect 17174 9068 17188 9082
rect 16637 9054 17188 9068
rect 16637 9052 16643 9054
rect 16614 9049 16643 9052
rect 16015 9034 16018 9040
rect 15932 9020 16018 9034
rect 16015 9014 16018 9020
rect 16044 9014 16047 9040
rect 17165 9014 17168 9040
rect 17194 9014 17197 9040
rect 19014 9034 19028 9083
rect 19290 9074 19304 9088
rect 19373 9082 19376 9108
rect 19402 9102 19405 9108
rect 19695 9102 19698 9108
rect 19402 9088 19698 9102
rect 19402 9082 19405 9088
rect 19695 9082 19698 9088
rect 19724 9102 19727 9108
rect 19834 9103 19863 9106
rect 19834 9102 19840 9103
rect 19724 9088 19840 9102
rect 19724 9082 19727 9088
rect 19834 9086 19840 9088
rect 19857 9086 19863 9103
rect 19834 9083 19863 9086
rect 19281 9048 19284 9074
rect 19310 9048 19313 9074
rect 20477 9034 20480 9040
rect 19014 9020 20480 9034
rect 20477 9014 20480 9020
rect 20506 9014 20509 9040
rect 20693 9034 20707 9122
rect 21995 9116 21998 9142
rect 22024 9136 22027 9142
rect 22602 9140 22616 9156
rect 22731 9150 22734 9156
rect 22760 9150 22763 9176
rect 23881 9150 23884 9176
rect 23910 9170 23913 9176
rect 24035 9171 24064 9174
rect 24035 9170 24041 9171
rect 23910 9156 24041 9170
rect 23910 9150 23913 9156
rect 24035 9154 24041 9156
rect 24058 9154 24064 9171
rect 24035 9151 24064 9154
rect 25675 9150 25678 9176
rect 25704 9170 25707 9176
rect 25859 9174 25862 9176
rect 25790 9171 25819 9174
rect 25790 9170 25796 9171
rect 25704 9156 25796 9170
rect 25704 9150 25707 9156
rect 25790 9154 25796 9156
rect 25813 9154 25819 9171
rect 25790 9151 25819 9154
rect 25841 9171 25862 9174
rect 25841 9154 25847 9171
rect 25841 9151 25862 9154
rect 25859 9150 25862 9151
rect 25888 9150 25891 9176
rect 26871 9150 26874 9176
rect 26900 9170 26903 9176
rect 26900 9156 27139 9170
rect 26900 9150 26903 9156
rect 22594 9137 22623 9140
rect 22594 9136 22600 9137
rect 22024 9122 22600 9136
rect 22024 9116 22027 9122
rect 22594 9120 22600 9122
rect 22617 9120 22623 9137
rect 22594 9117 22623 9120
rect 22639 9116 22642 9142
rect 22668 9136 22671 9142
rect 22686 9137 22715 9140
rect 22686 9136 22692 9137
rect 22668 9122 22692 9136
rect 22668 9116 22671 9122
rect 22686 9120 22692 9122
rect 22709 9120 22715 9137
rect 22686 9117 22715 9120
rect 22777 9116 22780 9142
rect 22806 9136 22809 9142
rect 23100 9137 23129 9140
rect 23100 9136 23106 9137
rect 22806 9122 23106 9136
rect 22806 9116 22809 9122
rect 23100 9120 23106 9122
rect 23123 9120 23129 9137
rect 23100 9117 23129 9120
rect 23330 9137 23359 9140
rect 23330 9120 23336 9137
rect 23353 9120 23359 9137
rect 23330 9117 23359 9120
rect 23338 9102 23352 9117
rect 23513 9116 23516 9142
rect 23542 9136 23545 9142
rect 23973 9136 23976 9142
rect 24002 9140 24005 9142
rect 24002 9137 24020 9140
rect 23542 9122 23976 9136
rect 23542 9116 23545 9122
rect 23973 9116 23976 9122
rect 24014 9120 24020 9137
rect 24002 9117 24020 9120
rect 24002 9116 24005 9117
rect 26917 9116 26920 9142
rect 26946 9116 26949 9142
rect 26975 9137 27004 9140
rect 26975 9136 26981 9137
rect 26972 9120 26981 9136
rect 26998 9120 27004 9137
rect 26972 9117 27004 9120
rect 22694 9088 23352 9102
rect 22694 9074 22708 9088
rect 23835 9082 23838 9108
rect 23864 9082 23867 9108
rect 25629 9082 25632 9108
rect 25658 9082 25661 9108
rect 26665 9103 26694 9106
rect 26665 9086 26671 9103
rect 26688 9102 26694 9103
rect 26972 9102 26986 9117
rect 27055 9116 27058 9142
rect 27084 9140 27087 9142
rect 27125 9140 27139 9156
rect 28021 9150 28024 9176
rect 28050 9170 28053 9176
rect 28274 9171 28303 9174
rect 28274 9170 28280 9171
rect 28050 9156 28280 9170
rect 28050 9150 28053 9156
rect 28274 9154 28280 9156
rect 28297 9154 28303 9171
rect 28274 9151 28303 9154
rect 28325 9171 28354 9174
rect 28325 9154 28331 9171
rect 28348 9170 28354 9171
rect 28348 9156 28458 9170
rect 28348 9154 28354 9156
rect 28325 9151 28354 9154
rect 28444 9142 28458 9156
rect 27239 9140 27242 9142
rect 27084 9137 27105 9140
rect 27099 9120 27105 9137
rect 27084 9117 27105 9120
rect 27124 9137 27153 9140
rect 27124 9120 27130 9137
rect 27147 9120 27153 9137
rect 27124 9117 27153 9120
rect 27179 9137 27208 9140
rect 27179 9120 27185 9137
rect 27202 9136 27208 9137
rect 27230 9137 27242 9140
rect 27202 9120 27216 9136
rect 27179 9117 27216 9120
rect 27230 9120 27236 9137
rect 27230 9117 27242 9120
rect 27084 9116 27087 9117
rect 26688 9088 26986 9102
rect 27202 9102 27216 9117
rect 27239 9116 27242 9117
rect 27268 9116 27271 9142
rect 27607 9116 27610 9142
rect 27636 9136 27639 9142
rect 27975 9136 27978 9142
rect 27636 9122 27978 9136
rect 27636 9116 27639 9122
rect 27975 9116 27978 9122
rect 28004 9136 28007 9142
rect 28114 9137 28143 9140
rect 28114 9136 28120 9137
rect 28004 9122 28120 9136
rect 28004 9116 28007 9122
rect 28114 9120 28120 9122
rect 28137 9120 28143 9137
rect 28114 9117 28143 9120
rect 28435 9116 28438 9142
rect 28464 9116 28467 9142
rect 27745 9102 27748 9108
rect 27202 9088 27748 9102
rect 26688 9086 26694 9088
rect 26665 9083 26694 9086
rect 27745 9082 27748 9088
rect 27774 9082 27777 9108
rect 22685 9048 22688 9074
rect 22714 9048 22717 9074
rect 24203 9034 24206 9040
rect 20693 9020 24206 9034
rect 24203 9014 24206 9020
rect 24232 9014 24235 9040
rect 25638 9034 25652 9082
rect 25813 9034 25816 9040
rect 25638 9020 25816 9034
rect 25813 9014 25816 9020
rect 25842 9014 25845 9040
rect 3036 8952 29992 9000
rect 14451 8912 14454 8938
rect 14480 8932 14483 8938
rect 14498 8933 14527 8936
rect 14498 8932 14504 8933
rect 14480 8918 14504 8932
rect 14480 8912 14483 8918
rect 14498 8916 14504 8918
rect 14521 8916 14527 8933
rect 14498 8913 14527 8916
rect 15969 8912 15972 8938
rect 15998 8912 16001 8938
rect 17855 8912 17858 8938
rect 17884 8912 17887 8938
rect 19925 8912 19928 8938
rect 19954 8932 19957 8938
rect 19954 8918 20546 8932
rect 19954 8912 19957 8918
rect 7782 8899 7811 8902
rect 7782 8882 7788 8899
rect 7805 8882 7811 8899
rect 7782 8879 7811 8882
rect 5896 8865 5925 8868
rect 5896 8848 5902 8865
rect 5919 8864 5925 8865
rect 5987 8864 5990 8870
rect 5919 8850 5990 8864
rect 5919 8848 5925 8850
rect 5896 8845 5925 8848
rect 5987 8844 5990 8850
rect 6016 8844 6019 8870
rect 6033 8844 6036 8870
rect 6062 8844 6065 8870
rect 7689 8844 7692 8870
rect 7718 8844 7721 8870
rect 7790 8864 7804 8879
rect 14129 8878 14132 8904
rect 14158 8898 14161 8904
rect 14405 8898 14408 8904
rect 14158 8884 14408 8898
rect 14158 8878 14161 8884
rect 14405 8878 14408 8884
rect 14434 8898 14437 8904
rect 20532 8898 20546 8918
rect 20707 8912 20710 8938
rect 20736 8936 20739 8938
rect 20736 8933 20760 8936
rect 20736 8916 20737 8933
rect 20754 8916 20760 8933
rect 27607 8932 27610 8938
rect 20736 8913 20760 8916
rect 26696 8918 27610 8932
rect 20736 8912 20739 8913
rect 22041 8898 22044 8904
rect 14434 8884 17947 8898
rect 20532 8884 22044 8898
rect 14434 8878 14437 8884
rect 7790 8850 8034 8864
rect 5619 8810 5622 8836
rect 5648 8830 5651 8836
rect 5850 8831 5879 8834
rect 5850 8830 5856 8831
rect 5648 8816 5856 8830
rect 5648 8810 5651 8816
rect 5850 8814 5856 8816
rect 5873 8830 5879 8831
rect 6079 8830 6082 8836
rect 5873 8816 6082 8830
rect 5873 8814 5879 8816
rect 5850 8811 5879 8814
rect 6079 8810 6082 8816
rect 6108 8810 6111 8836
rect 7598 8831 7627 8834
rect 7598 8814 7604 8831
rect 7621 8814 7627 8831
rect 7598 8811 7627 8814
rect 7782 8831 7811 8834
rect 7782 8814 7788 8831
rect 7805 8830 7811 8831
rect 7873 8830 7876 8836
rect 7805 8816 7876 8830
rect 7805 8814 7811 8816
rect 7782 8811 7811 8814
rect 7606 8796 7620 8811
rect 7873 8810 7876 8816
rect 7902 8810 7905 8836
rect 8020 8834 8034 8850
rect 9529 8844 9532 8870
rect 9558 8864 9561 8870
rect 10357 8864 10360 8870
rect 9558 8850 10360 8864
rect 9558 8844 9561 8850
rect 10357 8844 10360 8850
rect 10386 8844 10389 8870
rect 11093 8844 11096 8870
rect 11122 8864 11125 8870
rect 11370 8865 11399 8868
rect 11370 8864 11376 8865
rect 11122 8850 11376 8864
rect 11122 8844 11125 8850
rect 11370 8848 11376 8850
rect 11393 8848 11399 8865
rect 14590 8865 14619 8868
rect 14590 8864 14596 8865
rect 11370 8845 11399 8848
rect 14092 8850 14596 8864
rect 8012 8831 8041 8834
rect 8012 8814 8018 8831
rect 8035 8814 8041 8831
rect 8012 8811 8041 8814
rect 8103 8810 8106 8836
rect 8132 8810 8135 8836
rect 13440 8831 13469 8834
rect 13440 8814 13446 8831
rect 13463 8814 13469 8831
rect 13440 8811 13469 8814
rect 13574 8831 13603 8834
rect 13574 8814 13580 8831
rect 13597 8830 13603 8831
rect 14092 8830 14106 8850
rect 14590 8848 14596 8850
rect 14613 8848 14619 8865
rect 17933 8864 17947 8884
rect 22041 8878 22044 8884
rect 22070 8898 22073 8904
rect 22070 8884 25537 8898
rect 22070 8878 22073 8884
rect 18223 8864 18226 8870
rect 17933 8850 18226 8864
rect 14590 8845 14619 8848
rect 18223 8844 18226 8850
rect 18252 8844 18255 8870
rect 19695 8844 19698 8870
rect 19724 8844 19727 8870
rect 22639 8864 22642 8870
rect 22188 8850 22642 8864
rect 22188 8836 22202 8850
rect 22639 8844 22642 8850
rect 22668 8844 22671 8870
rect 13597 8816 14106 8830
rect 13597 8814 13603 8816
rect 13574 8811 13603 8814
rect 7827 8796 7830 8802
rect 7606 8782 7830 8796
rect 7827 8776 7830 8782
rect 7856 8776 7859 8802
rect 10496 8797 10525 8800
rect 10496 8780 10502 8797
rect 10519 8796 10525 8797
rect 10633 8796 10636 8802
rect 10519 8782 10636 8796
rect 10519 8780 10525 8782
rect 10496 8777 10525 8780
rect 10633 8776 10636 8782
rect 10662 8776 10665 8802
rect 10817 8776 10820 8802
rect 10846 8776 10849 8802
rect 11001 8776 11004 8802
rect 11030 8776 11033 8802
rect 13448 8796 13462 8811
rect 14313 8810 14316 8836
rect 14342 8830 14345 8836
rect 14406 8831 14435 8834
rect 14406 8830 14412 8831
rect 14342 8816 14412 8830
rect 14342 8810 14345 8816
rect 14406 8814 14412 8816
rect 14429 8814 14435 8831
rect 14406 8811 14435 8814
rect 14544 8831 14573 8834
rect 14544 8814 14550 8831
rect 14567 8814 14573 8831
rect 14544 8811 14573 8814
rect 13623 8796 13626 8802
rect 13448 8782 13626 8796
rect 13623 8776 13626 8782
rect 13652 8776 13655 8802
rect 13853 8776 13856 8802
rect 13882 8796 13885 8802
rect 14360 8797 14389 8800
rect 14360 8796 14366 8797
rect 13882 8782 14366 8796
rect 13882 8776 13885 8782
rect 14360 8780 14366 8782
rect 14383 8780 14389 8797
rect 14552 8796 14566 8811
rect 15095 8810 15098 8836
rect 15124 8830 15127 8836
rect 15124 8816 15762 8830
rect 15124 8810 15127 8816
rect 15233 8796 15236 8802
rect 14552 8782 15236 8796
rect 14360 8777 14389 8780
rect 15233 8776 15236 8782
rect 15262 8776 15265 8802
rect 15693 8776 15696 8802
rect 15722 8776 15725 8802
rect 15748 8796 15762 8816
rect 15785 8810 15788 8836
rect 15814 8810 15817 8836
rect 15831 8810 15834 8836
rect 15860 8810 15863 8836
rect 15878 8831 15907 8834
rect 15878 8814 15884 8831
rect 15901 8830 15907 8831
rect 17165 8830 17168 8836
rect 15901 8816 17168 8830
rect 15901 8814 15907 8816
rect 15878 8811 15907 8814
rect 17165 8810 17168 8816
rect 17194 8810 17197 8836
rect 17993 8810 17996 8836
rect 18022 8810 18025 8836
rect 19857 8831 19886 8834
rect 19857 8814 19863 8831
rect 19880 8830 19886 8831
rect 20109 8830 20112 8836
rect 19880 8816 20112 8830
rect 19880 8814 19886 8816
rect 19857 8811 19886 8814
rect 20109 8810 20112 8816
rect 20138 8810 20141 8836
rect 20247 8810 20250 8836
rect 20276 8830 20279 8836
rect 20385 8830 20388 8836
rect 20276 8816 20388 8830
rect 20276 8810 20279 8816
rect 20385 8810 20388 8816
rect 20414 8810 20417 8836
rect 22179 8810 22182 8836
rect 22208 8810 22211 8836
rect 22272 8831 22301 8834
rect 22272 8814 22278 8831
rect 22295 8814 22301 8831
rect 22272 8811 22301 8814
rect 22548 8831 22577 8834
rect 22548 8814 22554 8831
rect 22571 8830 22577 8831
rect 22777 8830 22780 8836
rect 22571 8816 22780 8830
rect 22571 8814 22577 8816
rect 22548 8811 22577 8814
rect 15970 8797 15999 8800
rect 15970 8796 15976 8797
rect 15748 8782 15976 8796
rect 15970 8780 15976 8782
rect 15993 8796 15999 8797
rect 16567 8796 16570 8802
rect 15993 8782 16570 8796
rect 15993 8780 15999 8782
rect 15970 8777 15999 8780
rect 16567 8776 16570 8782
rect 16596 8776 16599 8802
rect 17073 8776 17076 8802
rect 17102 8796 17105 8802
rect 17856 8797 17885 8800
rect 17856 8796 17862 8797
rect 17102 8782 17862 8796
rect 17102 8776 17105 8782
rect 17856 8780 17862 8782
rect 17879 8796 17885 8797
rect 19051 8796 19054 8802
rect 17879 8782 19054 8796
rect 17879 8780 17885 8782
rect 17856 8777 17885 8780
rect 19051 8776 19054 8782
rect 19080 8776 19083 8802
rect 19925 8800 19928 8802
rect 19907 8797 19928 8800
rect 19907 8780 19913 8797
rect 19907 8777 19928 8780
rect 19925 8776 19928 8777
rect 19954 8776 19957 8802
rect 21995 8776 21998 8802
rect 22024 8796 22027 8802
rect 22280 8796 22294 8811
rect 22777 8810 22780 8816
rect 22806 8810 22809 8836
rect 22824 8831 22853 8834
rect 22824 8814 22830 8831
rect 22847 8814 22853 8831
rect 25523 8830 25537 8884
rect 26696 8864 26710 8918
rect 27607 8912 27610 8918
rect 27636 8912 27639 8938
rect 27745 8912 27748 8938
rect 27774 8936 27777 8938
rect 27774 8933 27798 8936
rect 27774 8916 27775 8933
rect 27792 8916 27798 8933
rect 27774 8913 27798 8916
rect 27774 8912 27777 8913
rect 26734 8865 26763 8868
rect 26734 8864 26740 8865
rect 26696 8850 26740 8864
rect 26734 8848 26740 8850
rect 26757 8848 26763 8865
rect 26734 8845 26763 8848
rect 28343 8830 28346 8836
rect 25523 8816 28346 8830
rect 22824 8811 22853 8814
rect 22024 8782 22294 8796
rect 22024 8776 22027 8782
rect 22593 8776 22596 8802
rect 22622 8796 22625 8802
rect 22685 8796 22688 8802
rect 22622 8782 22688 8796
rect 22622 8776 22625 8782
rect 22685 8776 22688 8782
rect 22714 8796 22717 8802
rect 22832 8796 22846 8811
rect 22714 8782 22846 8796
rect 22714 8776 22717 8782
rect 25675 8776 25678 8802
rect 25704 8796 25707 8802
rect 26972 8800 26986 8816
rect 28343 8810 28346 8816
rect 28372 8810 28375 8836
rect 26895 8797 26924 8800
rect 26895 8796 26901 8797
rect 25704 8782 26901 8796
rect 25704 8776 25707 8782
rect 26895 8780 26901 8782
rect 26918 8780 26924 8797
rect 26895 8777 26924 8780
rect 26945 8797 26986 8800
rect 26945 8780 26951 8797
rect 26968 8782 26986 8797
rect 26968 8780 26974 8782
rect 26945 8777 26974 8780
rect 7643 8742 7646 8768
rect 7672 8742 7675 8768
rect 7781 8742 7784 8768
rect 7810 8762 7813 8768
rect 8058 8763 8087 8766
rect 8058 8762 8064 8763
rect 7810 8748 8064 8762
rect 7810 8742 7813 8748
rect 8058 8746 8064 8748
rect 8081 8746 8087 8763
rect 13632 8762 13646 8776
rect 14037 8762 14040 8768
rect 13632 8748 14040 8762
rect 8058 8743 8087 8746
rect 14037 8742 14040 8748
rect 14066 8742 14069 8768
rect 17948 8763 17977 8766
rect 17948 8746 17954 8763
rect 17971 8762 17977 8763
rect 18407 8762 18410 8768
rect 17971 8748 18410 8762
rect 17971 8746 17977 8748
rect 17948 8743 17977 8746
rect 18407 8742 18410 8748
rect 18436 8742 18439 8768
rect 22731 8742 22734 8768
rect 22760 8742 22763 8768
rect 23605 8742 23608 8768
rect 23634 8762 23637 8768
rect 25583 8762 25586 8768
rect 23634 8748 25586 8762
rect 23634 8742 23637 8748
rect 25583 8742 25586 8748
rect 25612 8742 25615 8768
rect 3036 8680 29992 8728
rect 7643 8640 7646 8666
rect 7672 8660 7675 8666
rect 7736 8661 7765 8664
rect 7736 8660 7742 8661
rect 7672 8646 7742 8660
rect 7672 8640 7675 8646
rect 7736 8644 7742 8646
rect 7759 8660 7765 8661
rect 7919 8660 7922 8666
rect 7759 8646 7922 8660
rect 7759 8644 7765 8646
rect 7736 8641 7765 8644
rect 7919 8640 7922 8646
rect 7948 8640 7951 8666
rect 9529 8640 9532 8666
rect 9558 8640 9561 8666
rect 10496 8661 10525 8664
rect 10496 8660 10502 8661
rect 10320 8646 10502 8660
rect 7827 8606 7830 8632
rect 7856 8606 7859 8632
rect 8012 8627 8041 8630
rect 8012 8610 8018 8627
rect 8035 8626 8041 8627
rect 8103 8626 8106 8632
rect 8035 8612 8106 8626
rect 8035 8610 8041 8612
rect 8012 8607 8041 8610
rect 8103 8606 8106 8612
rect 8132 8606 8135 8632
rect 8839 8606 8842 8632
rect 8868 8626 8871 8632
rect 9208 8627 9237 8630
rect 9208 8626 9214 8627
rect 8868 8612 9214 8626
rect 8868 8606 8871 8612
rect 9208 8610 9214 8612
rect 9231 8626 9237 8627
rect 10320 8626 10334 8646
rect 10496 8644 10502 8646
rect 10519 8660 10525 8661
rect 10519 8646 11024 8660
rect 10519 8644 10525 8646
rect 10496 8641 10525 8644
rect 9231 8612 10334 8626
rect 10458 8612 10610 8626
rect 9231 8610 9237 8612
rect 9208 8607 9237 8610
rect 10458 8598 10472 8612
rect 7735 8592 7738 8598
rect 7107 8578 7738 8592
rect 7735 8572 7738 8578
rect 7764 8572 7767 8598
rect 7782 8593 7811 8596
rect 7782 8576 7788 8593
rect 7805 8592 7811 8593
rect 7873 8592 7876 8598
rect 7805 8578 7876 8592
rect 7805 8576 7811 8578
rect 7782 8573 7811 8576
rect 7873 8572 7876 8578
rect 7902 8592 7905 8598
rect 8517 8592 8520 8598
rect 7902 8578 8520 8592
rect 7902 8572 7905 8578
rect 8517 8572 8520 8578
rect 8546 8592 8549 8598
rect 9070 8593 9099 8596
rect 9070 8592 9076 8593
rect 8546 8578 9076 8592
rect 8546 8572 8549 8578
rect 9070 8576 9076 8578
rect 9093 8576 9099 8593
rect 9070 8573 9099 8576
rect 9483 8572 9486 8598
rect 9512 8572 9515 8598
rect 10449 8572 10452 8598
rect 10478 8572 10481 8598
rect 10596 8592 10610 8612
rect 10633 8606 10636 8632
rect 10662 8626 10665 8632
rect 10680 8627 10709 8630
rect 10680 8626 10686 8627
rect 10662 8612 10686 8626
rect 10662 8606 10665 8612
rect 10680 8610 10686 8612
rect 10703 8610 10709 8627
rect 10680 8607 10709 8610
rect 11010 8596 11024 8646
rect 18407 8640 18410 8666
rect 18436 8640 18439 8666
rect 22869 8640 22872 8666
rect 22898 8640 22901 8666
rect 26849 8661 26878 8664
rect 26849 8644 26855 8661
rect 26872 8660 26878 8661
rect 27055 8660 27058 8666
rect 26872 8646 27058 8660
rect 26872 8644 26878 8646
rect 26849 8641 26878 8644
rect 27055 8640 27058 8646
rect 27084 8640 27087 8666
rect 21535 8606 21538 8632
rect 21564 8626 21567 8632
rect 23605 8630 23608 8632
rect 23583 8627 23608 8630
rect 23583 8626 23589 8627
rect 21564 8612 23589 8626
rect 21564 8606 21567 8612
rect 23583 8610 23589 8612
rect 23606 8610 23608 8627
rect 23583 8607 23608 8610
rect 23605 8606 23608 8607
rect 23634 8606 23637 8632
rect 25721 8606 25724 8632
rect 25750 8626 25753 8632
rect 26021 8627 26050 8630
rect 26021 8626 26027 8627
rect 25750 8612 26027 8626
rect 25750 8606 25753 8612
rect 26021 8610 26027 8612
rect 26044 8610 26050 8627
rect 26021 8607 26050 8610
rect 28803 8606 28806 8632
rect 28832 8606 28835 8632
rect 28850 8627 28879 8630
rect 28850 8610 28856 8627
rect 28873 8626 28879 8627
rect 28987 8626 28990 8632
rect 28873 8612 28990 8626
rect 28873 8610 28879 8612
rect 28850 8607 28879 8610
rect 28987 8606 28990 8612
rect 29016 8606 29019 8632
rect 10910 8593 10939 8596
rect 10910 8592 10916 8593
rect 10596 8578 10916 8592
rect 10910 8576 10916 8578
rect 10933 8576 10939 8593
rect 10910 8573 10939 8576
rect 11002 8593 11031 8596
rect 11002 8576 11008 8593
rect 11025 8592 11031 8593
rect 11047 8592 11050 8598
rect 11025 8578 11050 8592
rect 11025 8576 11031 8578
rect 11002 8573 11031 8576
rect 11047 8572 11050 8578
rect 11076 8572 11079 8598
rect 17073 8572 17076 8598
rect 17102 8572 17105 8598
rect 17165 8572 17168 8598
rect 17194 8572 17197 8598
rect 18223 8572 18226 8598
rect 18252 8592 18255 8598
rect 19235 8592 19238 8598
rect 18252 8578 19238 8592
rect 18252 8572 18255 8578
rect 19235 8572 19238 8578
rect 19264 8572 19267 8598
rect 21259 8572 21262 8598
rect 21288 8572 21291 8598
rect 21305 8572 21308 8598
rect 21334 8592 21337 8598
rect 21444 8593 21473 8596
rect 21444 8592 21450 8593
rect 21334 8578 21450 8592
rect 21334 8572 21337 8578
rect 21444 8576 21450 8578
rect 21467 8576 21473 8593
rect 21444 8573 21473 8576
rect 21627 8572 21630 8598
rect 21656 8572 21659 8598
rect 22042 8593 22071 8596
rect 22042 8576 22048 8593
rect 22065 8592 22071 8593
rect 22179 8592 22182 8598
rect 22065 8578 22182 8592
rect 22065 8576 22071 8578
rect 22042 8573 22071 8576
rect 22179 8572 22182 8578
rect 22208 8572 22211 8598
rect 22225 8572 22228 8598
rect 22254 8592 22257 8598
rect 22593 8592 22596 8598
rect 22254 8578 22596 8592
rect 22254 8572 22257 8578
rect 22593 8572 22596 8578
rect 22622 8572 22625 8598
rect 22639 8572 22642 8598
rect 22668 8592 22671 8598
rect 22732 8593 22761 8596
rect 22732 8592 22738 8593
rect 22668 8578 22738 8592
rect 22668 8572 22671 8578
rect 22732 8576 22738 8578
rect 22755 8576 22761 8593
rect 22732 8573 22761 8576
rect 22777 8572 22780 8598
rect 22806 8592 22809 8598
rect 22870 8593 22899 8596
rect 22870 8592 22876 8593
rect 22806 8578 22876 8592
rect 22806 8572 22809 8578
rect 22870 8576 22876 8578
rect 22893 8576 22899 8593
rect 22870 8573 22899 8576
rect 23237 8572 23240 8598
rect 23266 8592 23269 8598
rect 23376 8593 23405 8596
rect 23376 8592 23382 8593
rect 23266 8578 23382 8592
rect 23266 8572 23269 8578
rect 23376 8576 23382 8578
rect 23399 8576 23405 8593
rect 23376 8573 23405 8576
rect 23513 8572 23516 8598
rect 23542 8596 23545 8598
rect 23542 8593 23560 8596
rect 23554 8576 23560 8593
rect 23542 8573 23560 8576
rect 23542 8572 23545 8573
rect 25675 8572 25678 8598
rect 25704 8592 25707 8598
rect 25969 8593 25998 8596
rect 25969 8592 25975 8593
rect 25704 8578 25975 8592
rect 25704 8572 25707 8578
rect 25969 8576 25975 8578
rect 25992 8592 25998 8593
rect 28389 8592 28392 8598
rect 25992 8578 28392 8592
rect 25992 8576 25998 8578
rect 25969 8573 25998 8576
rect 28389 8572 28392 8578
rect 28418 8572 28421 8598
rect 28712 8593 28741 8596
rect 28712 8576 28718 8593
rect 28735 8576 28741 8593
rect 28712 8573 28741 8576
rect 6355 8538 6358 8564
rect 6384 8558 6387 8564
rect 6402 8559 6431 8562
rect 6402 8558 6408 8559
rect 6384 8544 6408 8558
rect 6384 8538 6387 8544
rect 6402 8542 6408 8544
rect 6425 8542 6431 8559
rect 6402 8539 6431 8542
rect 6539 8538 6542 8564
rect 6568 8538 6571 8564
rect 7414 8559 7443 8562
rect 7414 8542 7420 8559
rect 7437 8558 7443 8559
rect 7644 8559 7673 8562
rect 7644 8558 7650 8559
rect 7437 8544 7650 8558
rect 7437 8542 7443 8544
rect 7414 8539 7443 8542
rect 7644 8542 7650 8544
rect 7667 8558 7673 8559
rect 7689 8558 7692 8564
rect 7667 8544 7692 8558
rect 7667 8542 7673 8544
rect 7644 8539 7673 8542
rect 7689 8538 7692 8544
rect 7718 8538 7721 8564
rect 7744 8524 7758 8572
rect 8932 8559 8961 8562
rect 8932 8542 8938 8559
rect 8955 8558 8961 8559
rect 9115 8558 9118 8564
rect 8955 8544 9118 8558
rect 8955 8542 8961 8544
rect 8932 8539 8961 8542
rect 9115 8538 9118 8544
rect 9144 8538 9147 8564
rect 9162 8559 9191 8562
rect 9162 8542 9168 8559
rect 9185 8542 9191 8559
rect 9162 8539 9191 8542
rect 7873 8524 7876 8530
rect 7744 8510 7876 8524
rect 7873 8504 7876 8510
rect 7902 8504 7905 8530
rect 8885 8504 8888 8530
rect 8914 8524 8917 8530
rect 9024 8525 9053 8528
rect 9024 8524 9030 8525
rect 8914 8510 9030 8524
rect 8914 8504 8917 8510
rect 9024 8508 9030 8510
rect 9047 8508 9053 8525
rect 9024 8505 9053 8508
rect 8977 8470 8980 8496
rect 9006 8470 9009 8496
rect 9170 8490 9184 8539
rect 10633 8538 10636 8564
rect 10662 8538 10665 8564
rect 18269 8538 18272 8564
rect 18298 8538 18301 8564
rect 22961 8538 22964 8564
rect 22990 8538 22993 8564
rect 25813 8538 25816 8564
rect 25842 8538 25845 8564
rect 28720 8558 28734 8573
rect 28895 8572 28898 8598
rect 28924 8596 28927 8598
rect 28924 8592 28928 8596
rect 28924 8578 28946 8592
rect 28924 8573 28928 8578
rect 28924 8572 28927 8573
rect 29125 8558 29128 8564
rect 28720 8544 29128 8558
rect 29125 8538 29128 8544
rect 29154 8538 29157 8564
rect 10588 8525 10617 8528
rect 10588 8508 10594 8525
rect 10611 8524 10617 8525
rect 10910 8525 10939 8528
rect 10910 8524 10916 8525
rect 10611 8510 10916 8524
rect 10611 8508 10617 8510
rect 10588 8505 10617 8508
rect 10910 8508 10916 8510
rect 10933 8508 10939 8525
rect 10910 8505 10939 8508
rect 17119 8504 17122 8530
rect 17148 8524 17151 8530
rect 17212 8525 17241 8528
rect 17212 8524 17218 8525
rect 17148 8510 17218 8524
rect 17148 8504 17151 8510
rect 17212 8508 17218 8510
rect 17235 8508 17241 8525
rect 17212 8505 17241 8508
rect 21812 8525 21841 8528
rect 21812 8508 21818 8525
rect 21835 8524 21841 8525
rect 22133 8524 22136 8530
rect 21835 8510 22136 8524
rect 21835 8508 21841 8510
rect 21812 8505 21841 8508
rect 22133 8504 22136 8510
rect 22162 8504 22165 8530
rect 22685 8504 22688 8530
rect 22714 8524 22717 8530
rect 23100 8525 23129 8528
rect 23100 8524 23106 8525
rect 22714 8510 23106 8524
rect 22714 8504 22717 8510
rect 23100 8508 23106 8510
rect 23123 8508 23129 8525
rect 23100 8505 23129 8508
rect 27147 8504 27150 8530
rect 27176 8524 27179 8530
rect 28712 8525 28741 8528
rect 28712 8524 28718 8525
rect 27176 8510 28718 8524
rect 27176 8504 27179 8510
rect 28712 8508 28718 8510
rect 28735 8508 28741 8525
rect 28712 8505 28741 8508
rect 11093 8490 11096 8496
rect 9170 8476 11096 8490
rect 11093 8470 11096 8476
rect 11122 8470 11125 8496
rect 24341 8470 24344 8496
rect 24370 8490 24373 8496
rect 24411 8491 24440 8494
rect 24411 8490 24417 8491
rect 24370 8476 24417 8490
rect 24370 8470 24373 8476
rect 24411 8474 24417 8476
rect 24434 8474 24440 8491
rect 24411 8471 24440 8474
rect 3036 8408 29992 8456
rect 8517 8368 8520 8394
rect 8546 8368 8549 8394
rect 8932 8389 8961 8392
rect 8932 8372 8938 8389
rect 8955 8388 8961 8389
rect 9483 8388 9486 8394
rect 8955 8374 9486 8388
rect 8955 8372 8961 8374
rect 8932 8369 8961 8372
rect 9483 8368 9486 8374
rect 9512 8368 9515 8394
rect 24479 8388 24482 8394
rect 24442 8374 24482 8388
rect 19235 8334 19238 8360
rect 19264 8354 19267 8360
rect 20339 8354 20342 8360
rect 19264 8340 20342 8354
rect 19264 8334 19267 8340
rect 20339 8334 20342 8340
rect 20368 8354 20371 8360
rect 21259 8354 21262 8360
rect 20368 8340 21262 8354
rect 20368 8334 20371 8340
rect 21259 8334 21262 8340
rect 21288 8334 21291 8360
rect 24295 8334 24298 8360
rect 24324 8354 24327 8360
rect 24442 8354 24456 8374
rect 24479 8368 24482 8374
rect 24508 8388 24511 8394
rect 24508 8374 28987 8388
rect 24508 8368 24511 8374
rect 24324 8340 24456 8354
rect 24324 8334 24327 8340
rect 5850 8321 5879 8324
rect 5850 8304 5856 8321
rect 5873 8320 5879 8321
rect 6033 8320 6036 8326
rect 5873 8306 6036 8320
rect 5873 8304 5879 8306
rect 5850 8301 5879 8304
rect 6033 8300 6036 8306
rect 6062 8300 6065 8326
rect 6079 8300 6082 8326
rect 6108 8320 6111 8326
rect 6108 8306 6470 8320
rect 6108 8300 6111 8306
rect 5712 8287 5741 8290
rect 5712 8270 5718 8287
rect 5735 8270 5741 8287
rect 6456 8286 6470 8306
rect 7781 8300 7784 8326
rect 7810 8300 7813 8326
rect 20017 8300 20020 8326
rect 20046 8320 20049 8326
rect 20385 8320 20388 8326
rect 20046 8306 20388 8320
rect 20046 8300 20049 8306
rect 20385 8300 20388 8306
rect 20414 8300 20417 8326
rect 22142 8306 22616 8320
rect 6724 8287 6753 8290
rect 6724 8286 6730 8287
rect 6456 8272 6730 8286
rect 5712 8267 5741 8270
rect 6724 8270 6730 8272
rect 6747 8270 6753 8287
rect 6724 8267 6753 8270
rect 5720 8218 5734 8267
rect 7597 8266 7600 8292
rect 7626 8286 7629 8292
rect 7644 8287 7673 8290
rect 7644 8286 7650 8287
rect 7626 8272 7650 8286
rect 7626 8266 7629 8272
rect 7644 8270 7650 8272
rect 7667 8270 7673 8287
rect 7644 8267 7673 8270
rect 9392 8287 9421 8290
rect 9392 8270 9398 8287
rect 9415 8286 9421 8287
rect 9529 8286 9532 8292
rect 9415 8272 9532 8286
rect 9415 8270 9421 8272
rect 9392 8267 9421 8270
rect 9529 8266 9532 8272
rect 9558 8266 9561 8292
rect 19603 8266 19606 8292
rect 19632 8266 19635 8292
rect 19787 8266 19790 8292
rect 19816 8266 19819 8292
rect 19834 8287 19863 8290
rect 19834 8270 19840 8287
rect 19857 8270 19863 8287
rect 19834 8267 19863 8270
rect 19926 8287 19955 8290
rect 19926 8270 19932 8287
rect 19949 8286 19955 8287
rect 20891 8286 20894 8292
rect 19949 8272 20894 8286
rect 19949 8270 19955 8272
rect 19926 8267 19955 8270
rect 6079 8232 6082 8258
rect 6108 8232 6111 8258
rect 7882 8238 8027 8252
rect 7882 8224 7896 8238
rect 8747 8232 8750 8258
rect 8776 8252 8779 8258
rect 8794 8253 8823 8256
rect 8794 8252 8800 8253
rect 8776 8238 8800 8252
rect 8776 8232 8779 8238
rect 8794 8236 8800 8238
rect 8817 8236 8823 8253
rect 8794 8233 8823 8236
rect 19097 8232 19100 8258
rect 19126 8252 19129 8258
rect 19842 8252 19856 8267
rect 20891 8266 20894 8272
rect 20920 8266 20923 8292
rect 21305 8266 21308 8292
rect 21334 8286 21337 8292
rect 21995 8286 21998 8292
rect 21334 8272 21998 8286
rect 21334 8266 21337 8272
rect 21995 8266 21998 8272
rect 22024 8286 22027 8292
rect 22142 8290 22156 8306
rect 22134 8287 22163 8290
rect 22134 8286 22140 8287
rect 22024 8272 22140 8286
rect 22024 8266 22027 8272
rect 22134 8270 22140 8272
rect 22157 8270 22163 8287
rect 22134 8267 22163 8270
rect 22225 8266 22228 8292
rect 22254 8266 22257 8292
rect 22602 8286 22616 8306
rect 22639 8300 22642 8326
rect 22668 8320 22671 8326
rect 24442 8320 24456 8340
rect 22668 8306 22846 8320
rect 24442 8306 24485 8320
rect 22668 8300 22671 8306
rect 22685 8286 22688 8292
rect 22602 8272 22688 8286
rect 22685 8266 22688 8272
rect 22714 8266 22717 8292
rect 22732 8287 22761 8290
rect 22732 8270 22738 8287
rect 22755 8286 22761 8287
rect 22777 8286 22780 8292
rect 22755 8272 22780 8286
rect 22755 8270 22761 8272
rect 22732 8267 22761 8270
rect 22777 8266 22780 8272
rect 22806 8266 22809 8292
rect 22832 8286 22846 8306
rect 22870 8287 22899 8290
rect 22870 8286 22876 8287
rect 22832 8272 22876 8286
rect 22870 8270 22876 8272
rect 22893 8270 22899 8287
rect 22870 8267 22899 8270
rect 22961 8266 22964 8292
rect 22990 8286 22993 8292
rect 24341 8290 24344 8292
rect 24250 8287 24279 8290
rect 24250 8286 24256 8287
rect 22990 8272 24256 8286
rect 22990 8266 22993 8272
rect 24250 8270 24256 8272
rect 24273 8270 24279 8287
rect 24250 8267 24279 8270
rect 24327 8287 24344 8290
rect 24327 8270 24333 8287
rect 24327 8267 24344 8270
rect 24341 8266 24344 8267
rect 24370 8266 24373 8292
rect 24471 8290 24485 8306
rect 24387 8263 24390 8289
rect 24416 8288 24419 8289
rect 24416 8285 24430 8288
rect 24424 8268 24430 8285
rect 24416 8265 24430 8268
rect 24463 8287 24492 8290
rect 24463 8270 24469 8287
rect 24486 8270 24492 8287
rect 24463 8267 24492 8270
rect 24416 8263 24419 8265
rect 24510 8263 24513 8289
rect 24539 8263 24542 8289
rect 24562 8285 24591 8288
rect 24562 8268 24568 8285
rect 24585 8283 24591 8285
rect 24617 8283 24620 8292
rect 24585 8269 24620 8283
rect 24585 8268 24591 8269
rect 24562 8265 24591 8268
rect 24617 8266 24620 8269
rect 24646 8266 24649 8292
rect 28973 8286 28987 8374
rect 29355 8286 29358 8292
rect 28973 8272 29358 8286
rect 29355 8266 29358 8272
rect 29384 8266 29387 8292
rect 22915 8252 22918 8258
rect 19126 8238 19856 8252
rect 20693 8238 22918 8252
rect 19126 8232 19129 8238
rect 6355 8218 6358 8224
rect 5720 8204 6358 8218
rect 6355 8198 6358 8204
rect 6384 8218 6387 8224
rect 6861 8218 6864 8224
rect 6384 8204 6864 8218
rect 6384 8198 6387 8204
rect 6861 8198 6864 8204
rect 6890 8198 6893 8224
rect 7873 8198 7876 8224
rect 7902 8198 7905 8224
rect 8839 8198 8842 8224
rect 8868 8198 8871 8224
rect 20201 8198 20204 8224
rect 20230 8218 20233 8224
rect 20693 8218 20707 8238
rect 22915 8232 22918 8238
rect 22944 8232 22947 8258
rect 26825 8232 26828 8258
rect 26854 8252 26857 8258
rect 27377 8252 27380 8258
rect 26854 8238 27380 8252
rect 26854 8232 26857 8238
rect 27377 8232 27380 8238
rect 27406 8232 27409 8258
rect 20230 8204 20707 8218
rect 20230 8198 20233 8204
rect 22823 8198 22826 8224
rect 22852 8218 22855 8224
rect 22961 8218 22964 8224
rect 22852 8204 22964 8218
rect 22852 8198 22855 8204
rect 22961 8198 22964 8204
rect 22990 8198 22993 8224
rect 23007 8198 23010 8224
rect 23036 8218 23039 8224
rect 24295 8218 24298 8224
rect 23036 8204 24298 8218
rect 23036 8198 23039 8204
rect 24295 8198 24298 8204
rect 24324 8198 24327 8224
rect 24479 8198 24482 8224
rect 24508 8198 24511 8224
rect 3036 8136 29992 8184
rect 7689 8116 7692 8122
rect 6870 8102 7692 8116
rect 5987 8028 5990 8054
rect 6016 8048 6019 8054
rect 6402 8049 6431 8052
rect 6402 8048 6408 8049
rect 6016 8034 6408 8048
rect 6016 8028 6019 8034
rect 6402 8032 6408 8034
rect 6425 8032 6431 8049
rect 6402 8029 6431 8032
rect 6540 8049 6569 8052
rect 6540 8032 6546 8049
rect 6563 8048 6569 8049
rect 6585 8048 6588 8054
rect 6563 8034 6588 8048
rect 6563 8032 6569 8034
rect 6540 8029 6569 8032
rect 6585 8028 6588 8034
rect 6614 8028 6617 8054
rect 6632 8049 6661 8052
rect 6632 8032 6638 8049
rect 6655 8048 6661 8049
rect 6870 8048 6884 8102
rect 7689 8096 7692 8102
rect 7718 8096 7721 8122
rect 7873 8116 7876 8122
rect 7744 8102 7876 8116
rect 7744 8088 7758 8102
rect 7873 8096 7876 8102
rect 7902 8096 7905 8122
rect 15510 8117 15539 8120
rect 15510 8100 15516 8117
rect 15533 8116 15539 8117
rect 15693 8116 15696 8122
rect 15533 8102 15696 8116
rect 15533 8100 15539 8102
rect 15510 8097 15539 8100
rect 15693 8096 15696 8102
rect 15722 8096 15725 8122
rect 17350 8117 17379 8120
rect 17350 8100 17356 8117
rect 17373 8116 17379 8117
rect 17993 8116 17996 8122
rect 17373 8102 17996 8116
rect 17373 8100 17379 8102
rect 17350 8097 17379 8100
rect 17993 8096 17996 8102
rect 18022 8096 18025 8122
rect 18269 8096 18272 8122
rect 18298 8116 18301 8122
rect 18592 8117 18621 8120
rect 18592 8116 18598 8117
rect 18298 8102 18598 8116
rect 18298 8096 18301 8102
rect 18592 8100 18598 8102
rect 18615 8100 18621 8117
rect 18592 8097 18621 8100
rect 19281 8096 19284 8122
rect 19310 8116 19313 8122
rect 21029 8116 21032 8122
rect 19310 8102 20408 8116
rect 19310 8096 19313 8102
rect 7735 8082 7738 8088
rect 7613 8068 7738 8082
rect 7735 8062 7738 8068
rect 7764 8062 7767 8088
rect 7827 8062 7830 8088
rect 7856 8082 7859 8088
rect 20156 8083 20185 8086
rect 7856 8068 8264 8082
rect 7856 8062 7859 8068
rect 8104 8049 8133 8052
rect 8104 8048 8110 8049
rect 6655 8034 6884 8048
rect 7928 8034 8110 8048
rect 6655 8032 6661 8034
rect 6632 8029 6661 8032
rect 7928 8020 7942 8034
rect 8104 8032 8110 8034
rect 8127 8032 8133 8049
rect 8104 8029 8133 8032
rect 8195 8028 8198 8054
rect 8224 8028 8227 8054
rect 8250 8052 8264 8068
rect 20156 8066 20162 8083
rect 20179 8082 20185 8083
rect 20201 8082 20204 8088
rect 20179 8068 20204 8082
rect 20179 8066 20185 8068
rect 20156 8063 20185 8066
rect 20201 8062 20204 8068
rect 20230 8062 20233 8088
rect 20394 8086 20408 8102
rect 20624 8102 21032 8116
rect 20386 8083 20415 8086
rect 20386 8066 20392 8083
rect 20409 8066 20415 8083
rect 20386 8063 20415 8066
rect 8242 8049 8271 8052
rect 8242 8032 8248 8049
rect 8265 8032 8271 8049
rect 8242 8029 8271 8032
rect 10449 8028 10452 8054
rect 10478 8048 10481 8054
rect 10587 8048 10590 8054
rect 10478 8034 10590 8048
rect 10478 8028 10481 8034
rect 10587 8028 10590 8034
rect 10616 8048 10619 8054
rect 10726 8049 10755 8052
rect 10726 8048 10732 8049
rect 10616 8034 10732 8048
rect 10616 8028 10619 8034
rect 10726 8032 10732 8034
rect 10749 8032 10755 8049
rect 10726 8029 10755 8032
rect 14405 8028 14408 8054
rect 14434 8028 14437 8054
rect 14497 8028 14500 8054
rect 14526 8028 14529 8054
rect 14543 8028 14546 8054
rect 14572 8028 14575 8054
rect 15326 8049 15355 8052
rect 15326 8032 15332 8049
rect 15349 8048 15355 8049
rect 16107 8048 16110 8054
rect 15349 8034 16110 8048
rect 15349 8032 15355 8034
rect 15326 8029 15355 8032
rect 16107 8028 16110 8034
rect 16136 8028 16139 8054
rect 17166 8049 17195 8052
rect 17166 8032 17172 8049
rect 17189 8048 17195 8049
rect 17487 8048 17490 8054
rect 17189 8034 17490 8048
rect 17189 8032 17195 8034
rect 17166 8029 17195 8032
rect 17487 8028 17490 8034
rect 17516 8028 17519 8054
rect 18085 8028 18088 8054
rect 18114 8048 18117 8054
rect 18408 8049 18437 8052
rect 18408 8048 18414 8049
rect 18114 8034 18414 8048
rect 18114 8028 18117 8034
rect 18408 8032 18414 8034
rect 18431 8032 18437 8049
rect 18408 8029 18437 8032
rect 18637 8028 18640 8054
rect 18666 8048 18669 8054
rect 20110 8049 20139 8052
rect 20110 8048 20116 8049
rect 18666 8034 20116 8048
rect 18666 8028 18669 8034
rect 20110 8032 20116 8034
rect 20133 8032 20139 8049
rect 20110 8029 20139 8032
rect 6861 7994 6864 8020
rect 6890 7994 6893 8020
rect 7000 8015 7029 8018
rect 7000 7998 7006 8015
rect 7023 8014 7029 8015
rect 7643 8014 7646 8020
rect 7023 8000 7646 8014
rect 7023 7998 7029 8000
rect 7000 7995 7029 7998
rect 7643 7994 7646 8000
rect 7672 7994 7675 8020
rect 7689 7994 7692 8020
rect 7718 7994 7721 8020
rect 7874 8015 7903 8018
rect 7874 7998 7880 8015
rect 7897 8014 7903 8015
rect 7919 8014 7922 8020
rect 7897 8000 7922 8014
rect 7897 7998 7903 8000
rect 7874 7995 7903 7998
rect 7919 7994 7922 8000
rect 7948 7994 7951 8020
rect 10403 7994 10406 8020
rect 10432 8014 10435 8020
rect 10633 8014 10636 8020
rect 10432 8000 10636 8014
rect 10432 7994 10435 8000
rect 10633 7994 10636 8000
rect 10662 8014 10665 8020
rect 10864 8015 10893 8018
rect 10864 8014 10870 8015
rect 10662 8000 10870 8014
rect 10662 7994 10665 8000
rect 10864 7998 10870 8000
rect 10887 7998 10893 8015
rect 10864 7995 10893 7998
rect 13853 7994 13856 8020
rect 13882 8014 13885 8020
rect 15280 8015 15309 8018
rect 15280 8014 15286 8015
rect 13882 8000 15286 8014
rect 13882 7994 13885 8000
rect 15280 7998 15286 8000
rect 15303 7998 15309 8015
rect 15280 7995 15309 7998
rect 15877 7994 15880 8020
rect 15906 8014 15909 8020
rect 15969 8014 15972 8020
rect 15906 8000 15972 8014
rect 15906 7994 15909 8000
rect 15969 7994 15972 8000
rect 15998 8014 16001 8020
rect 17120 8015 17149 8018
rect 17120 8014 17126 8015
rect 15998 8000 17126 8014
rect 15998 7994 16001 8000
rect 17120 7998 17126 8000
rect 17143 7998 17149 8015
rect 17120 7995 17149 7998
rect 17395 7994 17398 8020
rect 17424 7994 17427 8020
rect 18454 8015 18483 8018
rect 18454 7998 18460 8015
rect 18477 8014 18483 8015
rect 19327 8014 19330 8020
rect 18477 8000 19330 8014
rect 18477 7998 18483 8000
rect 18454 7995 18483 7998
rect 19327 7994 19330 8000
rect 19356 7994 19359 8020
rect 6402 7981 6431 7984
rect 6402 7964 6408 7981
rect 6425 7980 6431 7981
rect 7698 7980 7712 7994
rect 8195 7980 8198 7986
rect 6425 7966 6930 7980
rect 7698 7966 8198 7980
rect 6425 7964 6431 7966
rect 6402 7961 6431 7964
rect 6540 7947 6569 7950
rect 6540 7930 6546 7947
rect 6563 7946 6569 7947
rect 6815 7946 6818 7952
rect 6563 7932 6818 7946
rect 6563 7930 6569 7932
rect 6540 7927 6569 7930
rect 6815 7926 6818 7932
rect 6844 7926 6847 7952
rect 6916 7946 6930 7966
rect 8195 7960 8198 7966
rect 8224 7960 8227 7986
rect 10772 7981 10801 7984
rect 10772 7964 10778 7981
rect 10795 7980 10801 7981
rect 11553 7980 11556 7986
rect 10795 7966 11556 7980
rect 10795 7964 10801 7966
rect 10772 7961 10801 7964
rect 11553 7960 11556 7966
rect 11582 7960 11585 7986
rect 17165 7960 17168 7986
rect 17194 7980 17197 7986
rect 17350 7981 17379 7984
rect 17350 7980 17356 7981
rect 17194 7966 17356 7980
rect 17194 7960 17197 7966
rect 17350 7964 17356 7966
rect 17373 7964 17379 7981
rect 20118 7980 20132 8029
rect 20339 8028 20342 8054
rect 20368 8028 20371 8054
rect 20394 8048 20408 8063
rect 20431 8062 20434 8088
rect 20460 8082 20463 8088
rect 20624 8082 20638 8102
rect 21029 8096 21032 8102
rect 21058 8116 21061 8122
rect 21305 8116 21308 8122
rect 21058 8102 21308 8116
rect 21058 8096 21061 8102
rect 20460 8068 20638 8082
rect 20693 8068 21098 8082
rect 20460 8062 20463 8068
rect 20693 8048 20707 8068
rect 21084 8054 21098 8068
rect 20394 8034 20707 8048
rect 20753 8028 20756 8054
rect 20782 8048 20785 8054
rect 20800 8049 20829 8052
rect 20800 8048 20806 8049
rect 20782 8034 20806 8048
rect 20782 8028 20785 8034
rect 20800 8032 20806 8034
rect 20823 8032 20829 8049
rect 20800 8029 20829 8032
rect 21075 8028 21078 8054
rect 21104 8028 21107 8054
rect 21176 8052 21190 8102
rect 21305 8096 21308 8102
rect 21334 8096 21337 8122
rect 21351 8096 21354 8122
rect 21380 8096 21383 8122
rect 22731 8096 22734 8122
rect 22760 8116 22763 8122
rect 23007 8116 23010 8122
rect 22760 8102 23010 8116
rect 22760 8096 22763 8102
rect 23007 8096 23010 8102
rect 23036 8096 23039 8122
rect 24227 8117 24256 8120
rect 24227 8100 24233 8117
rect 24250 8116 24256 8117
rect 24387 8116 24390 8122
rect 24250 8102 24390 8116
rect 24250 8100 24256 8102
rect 24227 8097 24256 8100
rect 24387 8096 24390 8102
rect 24416 8096 24419 8122
rect 24479 8096 24482 8122
rect 24508 8116 24511 8122
rect 24756 8117 24785 8120
rect 24756 8116 24762 8117
rect 24508 8102 24762 8116
rect 24508 8096 24511 8102
rect 24756 8100 24762 8102
rect 24779 8100 24785 8117
rect 24756 8097 24785 8100
rect 24801 8096 24804 8122
rect 24830 8096 24833 8122
rect 29125 8096 29128 8122
rect 29154 8120 29157 8122
rect 29154 8117 29178 8120
rect 29154 8100 29155 8117
rect 29172 8100 29178 8117
rect 29154 8097 29178 8100
rect 29154 8096 29157 8097
rect 23421 8086 23424 8088
rect 23403 8083 23424 8086
rect 23403 8066 23409 8083
rect 23403 8063 23424 8066
rect 23421 8062 23424 8063
rect 23450 8062 23453 8088
rect 28343 8086 28346 8088
rect 28325 8083 28346 8086
rect 28325 8066 28331 8083
rect 28325 8063 28346 8066
rect 28343 8062 28346 8063
rect 28372 8062 28375 8088
rect 21168 8049 21197 8052
rect 21168 8032 21174 8049
rect 21191 8032 21197 8049
rect 21168 8029 21197 8032
rect 21536 8049 21565 8052
rect 21536 8032 21542 8049
rect 21559 8048 21565 8049
rect 21627 8048 21630 8054
rect 21559 8034 21630 8048
rect 21559 8032 21565 8034
rect 21536 8029 21565 8032
rect 20348 8014 20362 8028
rect 20762 8014 20776 8028
rect 21544 8014 21558 8029
rect 21627 8028 21630 8034
rect 21656 8028 21659 8054
rect 23192 8049 23221 8052
rect 23192 8032 23198 8049
rect 23215 8048 23221 8049
rect 23237 8048 23240 8054
rect 23215 8034 23240 8048
rect 23215 8032 23221 8034
rect 23192 8029 23221 8032
rect 23237 8028 23240 8034
rect 23266 8028 23269 8054
rect 23353 8049 23382 8052
rect 23353 8032 23359 8049
rect 23376 8048 23382 8049
rect 23513 8048 23516 8054
rect 23376 8034 23516 8048
rect 23376 8032 23382 8034
rect 23353 8029 23382 8032
rect 23513 8028 23516 8034
rect 23542 8028 23545 8054
rect 24709 8028 24712 8054
rect 24738 8028 24741 8054
rect 24894 8049 24923 8052
rect 24894 8032 24900 8049
rect 24917 8048 24923 8049
rect 25261 8048 25264 8054
rect 24917 8034 25264 8048
rect 24917 8032 24923 8034
rect 24894 8029 24923 8032
rect 25261 8028 25264 8034
rect 25290 8028 25293 8054
rect 28067 8028 28070 8054
rect 28096 8048 28099 8054
rect 28275 8049 28304 8052
rect 28275 8048 28281 8049
rect 28096 8034 28281 8048
rect 28096 8028 28099 8034
rect 28275 8032 28281 8034
rect 28298 8048 28304 8049
rect 28389 8048 28392 8054
rect 28298 8034 28392 8048
rect 28298 8032 28304 8034
rect 28275 8029 28304 8032
rect 28389 8028 28392 8034
rect 28418 8028 28421 8054
rect 20348 8000 20776 8014
rect 20992 8000 21558 8014
rect 20992 7986 21006 8000
rect 22133 7994 22136 8020
rect 22162 8014 22165 8020
rect 22271 8014 22274 8020
rect 22162 8000 22274 8014
rect 22162 7994 22165 8000
rect 22271 7994 22274 8000
rect 22300 7994 22303 8020
rect 27975 7994 27978 8020
rect 28004 8014 28007 8020
rect 28114 8015 28143 8018
rect 28114 8014 28120 8015
rect 28004 8000 28120 8014
rect 28004 7994 28007 8000
rect 28114 7998 28120 8000
rect 28137 7998 28143 8015
rect 28114 7995 28143 7998
rect 20983 7980 20986 7986
rect 20118 7966 20986 7980
rect 17350 7961 17379 7964
rect 20983 7960 20986 7966
rect 21012 7960 21015 7986
rect 24755 7960 24758 7986
rect 24784 7960 24787 7986
rect 7689 7946 7692 7952
rect 6916 7932 7692 7946
rect 7689 7926 7692 7932
rect 7718 7926 7721 7952
rect 8103 7926 8106 7952
rect 8132 7926 8135 7952
rect 10679 7926 10682 7952
rect 10708 7946 10711 7952
rect 10726 7947 10755 7950
rect 10726 7946 10732 7947
rect 10708 7932 10732 7946
rect 10708 7926 10711 7932
rect 10726 7930 10732 7932
rect 10749 7930 10755 7947
rect 10726 7927 10755 7930
rect 13715 7926 13718 7952
rect 13744 7946 13747 7952
rect 14314 7947 14343 7950
rect 14314 7946 14320 7947
rect 13744 7932 14320 7946
rect 13744 7926 13747 7932
rect 14314 7930 14320 7932
rect 14337 7930 14343 7947
rect 14314 7927 14343 7930
rect 20753 7926 20756 7952
rect 20782 7946 20785 7952
rect 22133 7946 22136 7952
rect 20782 7932 22136 7946
rect 20782 7926 20785 7932
rect 22133 7926 22136 7932
rect 22162 7946 22165 7952
rect 22225 7946 22228 7952
rect 22162 7932 22228 7946
rect 22162 7926 22165 7932
rect 22225 7926 22228 7932
rect 22254 7926 22257 7952
rect 3036 7864 29992 7912
rect 6539 7824 6542 7850
rect 6568 7844 6571 7850
rect 6816 7845 6845 7848
rect 6816 7844 6822 7845
rect 6568 7830 6822 7844
rect 6568 7824 6571 7830
rect 6816 7828 6822 7830
rect 6839 7828 6845 7845
rect 6816 7825 6845 7828
rect 7598 7845 7627 7848
rect 7598 7828 7604 7845
rect 7621 7844 7627 7845
rect 8103 7844 8106 7850
rect 7621 7830 8106 7844
rect 7621 7828 7627 7830
rect 7598 7825 7627 7828
rect 8103 7824 8106 7830
rect 8132 7824 8135 7850
rect 15969 7824 15972 7850
rect 15998 7824 16001 7850
rect 17487 7824 17490 7850
rect 17516 7824 17519 7850
rect 19649 7824 19652 7850
rect 19678 7844 19681 7850
rect 28343 7844 28346 7850
rect 19678 7830 28346 7844
rect 19678 7824 19681 7830
rect 28343 7824 28346 7830
rect 28372 7824 28375 7850
rect 28987 7848 28990 7850
rect 28965 7845 28990 7848
rect 28965 7828 28971 7845
rect 28988 7828 28990 7845
rect 28965 7825 28990 7828
rect 28987 7824 28990 7825
rect 29016 7824 29019 7850
rect 29033 7824 29036 7850
rect 29062 7844 29065 7850
rect 29494 7845 29523 7848
rect 29494 7844 29500 7845
rect 29062 7830 29500 7844
rect 29062 7824 29065 7830
rect 29494 7828 29500 7830
rect 29517 7828 29523 7845
rect 29494 7825 29523 7828
rect 7643 7790 7646 7816
rect 7672 7790 7675 7816
rect 14497 7790 14500 7816
rect 14526 7810 14529 7816
rect 19281 7810 19284 7816
rect 14526 7796 19284 7810
rect 14526 7790 14529 7796
rect 6585 7756 6588 7782
rect 6614 7776 6617 7782
rect 7781 7776 7784 7782
rect 6614 7762 6976 7776
rect 6614 7756 6617 7762
rect 6815 7722 6818 7748
rect 6844 7722 6847 7748
rect 6962 7746 6976 7762
rect 7422 7762 7784 7776
rect 7422 7746 7436 7762
rect 7781 7756 7784 7762
rect 7810 7756 7813 7782
rect 10357 7756 10360 7782
rect 10386 7776 10389 7782
rect 10542 7777 10571 7780
rect 10542 7776 10548 7777
rect 10386 7762 10548 7776
rect 10386 7756 10389 7762
rect 10542 7760 10548 7762
rect 10565 7760 10571 7777
rect 10542 7757 10571 7760
rect 10679 7756 10682 7782
rect 10708 7756 10711 7782
rect 14037 7776 14040 7782
rect 13816 7762 14040 7776
rect 6954 7743 6983 7746
rect 6954 7726 6960 7743
rect 6977 7742 6983 7743
rect 7414 7743 7443 7746
rect 7414 7742 7420 7743
rect 6977 7728 7420 7742
rect 6977 7726 6983 7728
rect 6954 7723 6983 7726
rect 7414 7726 7420 7728
rect 7437 7726 7443 7743
rect 7414 7723 7443 7726
rect 7644 7743 7673 7746
rect 7644 7726 7650 7743
rect 7667 7742 7673 7743
rect 7689 7742 7692 7748
rect 7667 7728 7692 7742
rect 7667 7726 7673 7728
rect 7644 7723 7673 7726
rect 7689 7722 7692 7728
rect 7718 7742 7721 7748
rect 10403 7742 10406 7748
rect 7718 7728 10406 7742
rect 7718 7722 7721 7728
rect 10403 7722 10406 7728
rect 10432 7722 10435 7748
rect 13715 7722 13718 7748
rect 13744 7722 13747 7748
rect 13816 7746 13830 7762
rect 14037 7756 14040 7762
rect 14066 7776 14069 7782
rect 14130 7777 14159 7780
rect 14130 7776 14136 7777
rect 14066 7762 14136 7776
rect 14066 7756 14069 7762
rect 14130 7760 14136 7762
rect 14153 7760 14159 7777
rect 14506 7776 14520 7790
rect 14130 7757 14159 7760
rect 14276 7762 14520 7776
rect 15740 7777 15769 7780
rect 13808 7743 13837 7746
rect 13808 7726 13814 7743
rect 13831 7726 13837 7743
rect 13808 7723 13837 7726
rect 13853 7722 13856 7748
rect 13882 7722 13885 7748
rect 14276 7746 14290 7762
rect 15740 7760 15746 7777
rect 15763 7760 15769 7777
rect 15740 7757 15769 7760
rect 14084 7743 14113 7746
rect 14084 7726 14090 7743
rect 14107 7726 14113 7743
rect 14084 7723 14113 7726
rect 14268 7743 14297 7746
rect 14268 7726 14274 7743
rect 14291 7726 14297 7743
rect 14268 7723 14297 7726
rect 14360 7743 14389 7746
rect 14360 7726 14366 7743
rect 14383 7742 14389 7743
rect 14543 7742 14546 7748
rect 14383 7728 14546 7742
rect 14383 7726 14389 7728
rect 14360 7723 14389 7726
rect 7460 7709 7489 7712
rect 7460 7692 7466 7709
rect 7483 7708 7489 7709
rect 7919 7708 7922 7714
rect 7483 7694 7922 7708
rect 7483 7692 7489 7694
rect 7460 7689 7489 7692
rect 7919 7688 7922 7694
rect 7948 7688 7951 7714
rect 11001 7688 11004 7714
rect 11030 7688 11033 7714
rect 11507 7688 11510 7714
rect 11536 7708 11539 7714
rect 11554 7709 11583 7712
rect 11554 7708 11560 7709
rect 11536 7694 11560 7708
rect 11536 7688 11539 7694
rect 11554 7692 11560 7694
rect 11577 7692 11583 7709
rect 14092 7708 14106 7723
rect 14543 7722 14546 7728
rect 14572 7742 14575 7748
rect 15748 7742 15762 7757
rect 14572 7728 15762 7742
rect 15786 7743 15815 7746
rect 14572 7722 14575 7728
rect 15786 7726 15792 7743
rect 15809 7742 15815 7743
rect 15969 7742 15972 7748
rect 15809 7728 15972 7742
rect 15809 7726 15815 7728
rect 15786 7723 15815 7726
rect 15969 7722 15972 7728
rect 15998 7722 16001 7748
rect 17358 7746 17372 7796
rect 19281 7790 19284 7796
rect 19310 7790 19313 7816
rect 20017 7790 20020 7816
rect 20046 7810 20049 7816
rect 20201 7810 20204 7816
rect 20046 7796 20204 7810
rect 20046 7790 20049 7796
rect 20201 7790 20204 7796
rect 20230 7810 20233 7816
rect 20230 7796 21236 7810
rect 20230 7790 20233 7796
rect 17396 7777 17425 7780
rect 17396 7760 17402 7777
rect 17419 7776 17425 7777
rect 18269 7776 18272 7782
rect 17419 7762 18272 7776
rect 17419 7760 17425 7762
rect 17396 7757 17425 7760
rect 18269 7756 18272 7762
rect 18298 7756 18301 7782
rect 19420 7777 19449 7780
rect 19060 7762 19350 7776
rect 17350 7743 17379 7746
rect 17350 7726 17356 7743
rect 17373 7726 17379 7743
rect 17350 7723 17379 7726
rect 18315 7722 18318 7748
rect 18344 7742 18347 7748
rect 19060 7746 19074 7762
rect 19052 7743 19081 7746
rect 19052 7742 19058 7743
rect 18344 7728 19058 7742
rect 18344 7722 18347 7728
rect 19052 7726 19058 7728
rect 19075 7726 19081 7743
rect 19052 7723 19081 7726
rect 19143 7722 19146 7748
rect 19172 7742 19175 7748
rect 19282 7743 19311 7746
rect 19282 7742 19288 7743
rect 19172 7728 19288 7742
rect 19172 7722 19175 7728
rect 19282 7726 19288 7728
rect 19305 7726 19311 7743
rect 19336 7742 19350 7762
rect 19420 7760 19426 7777
rect 19443 7776 19449 7777
rect 20937 7776 20940 7782
rect 19443 7762 20940 7776
rect 19443 7760 19449 7762
rect 19420 7757 19449 7760
rect 20937 7756 20940 7762
rect 20966 7756 20969 7782
rect 19972 7743 20001 7746
rect 19972 7742 19978 7743
rect 19336 7728 19978 7742
rect 19282 7723 19311 7726
rect 19972 7726 19978 7728
rect 19995 7742 20001 7743
rect 20017 7742 20020 7748
rect 19995 7728 20020 7742
rect 19995 7726 20001 7728
rect 19972 7723 20001 7726
rect 20017 7722 20020 7728
rect 20046 7722 20049 7748
rect 21222 7746 21236 7796
rect 22271 7790 22274 7816
rect 22300 7810 22303 7816
rect 22300 7796 23214 7810
rect 22300 7790 22303 7796
rect 21535 7756 21538 7782
rect 21564 7756 21567 7782
rect 21627 7756 21630 7782
rect 21656 7776 21659 7782
rect 22777 7776 22780 7782
rect 21656 7762 22780 7776
rect 21656 7756 21659 7762
rect 20110 7743 20139 7746
rect 20110 7726 20116 7743
rect 20133 7726 20139 7743
rect 20110 7723 20139 7726
rect 21214 7743 21243 7746
rect 21214 7726 21220 7743
rect 21237 7726 21243 7743
rect 21214 7723 21243 7726
rect 14405 7708 14408 7714
rect 14092 7694 14408 7708
rect 11554 7689 11583 7692
rect 14405 7688 14408 7694
rect 14434 7688 14437 7714
rect 19097 7688 19100 7714
rect 19126 7708 19129 7714
rect 20118 7708 20132 7723
rect 21443 7722 21446 7748
rect 21472 7722 21475 7748
rect 22088 7743 22117 7746
rect 22088 7726 22094 7743
rect 22111 7742 22117 7743
rect 22133 7742 22136 7748
rect 22111 7728 22136 7742
rect 22111 7726 22117 7728
rect 22088 7723 22117 7726
rect 22133 7722 22136 7728
rect 22162 7722 22165 7748
rect 22179 7722 22182 7748
rect 22208 7722 22211 7748
rect 22602 7746 22616 7762
rect 22777 7756 22780 7762
rect 22806 7756 22809 7782
rect 23200 7776 23214 7796
rect 24801 7790 24804 7816
rect 24830 7810 24833 7816
rect 26734 7811 26763 7814
rect 26734 7810 26740 7811
rect 24830 7796 26740 7810
rect 24830 7790 24833 7796
rect 26734 7794 26740 7796
rect 26757 7794 26763 7811
rect 26734 7791 26763 7794
rect 23200 7762 24157 7776
rect 22594 7743 22623 7746
rect 22594 7726 22600 7743
rect 22617 7726 22623 7743
rect 22594 7723 22623 7726
rect 22685 7722 22688 7748
rect 22714 7742 22717 7748
rect 22824 7743 22853 7746
rect 22824 7742 22830 7743
rect 22714 7728 22830 7742
rect 22714 7722 22717 7728
rect 22824 7726 22830 7728
rect 22847 7726 22853 7743
rect 22824 7723 22853 7726
rect 19126 7694 20132 7708
rect 19126 7688 19129 7694
rect 21075 7688 21078 7714
rect 21104 7708 21107 7714
rect 22188 7708 22202 7722
rect 21104 7694 22202 7708
rect 24143 7708 24157 7762
rect 26733 7722 26736 7748
rect 26762 7722 26765 7748
rect 26825 7746 26828 7748
rect 26811 7743 26828 7746
rect 26811 7726 26817 7743
rect 26811 7723 26828 7726
rect 26825 7722 26828 7723
rect 26854 7722 26857 7748
rect 26995 7743 27024 7746
rect 26895 7733 26924 7736
rect 26895 7716 26901 7733
rect 26918 7716 26924 7733
rect 26895 7714 26924 7716
rect 24143 7694 26833 7708
rect 21104 7688 21107 7694
rect 6908 7675 6937 7678
rect 6908 7658 6914 7675
rect 6931 7674 6937 7675
rect 7506 7675 7535 7678
rect 7506 7674 7512 7675
rect 6931 7660 7512 7674
rect 6931 7658 6937 7660
rect 6908 7655 6937 7658
rect 7506 7658 7512 7660
rect 7529 7674 7535 7675
rect 7827 7674 7830 7680
rect 7529 7660 7830 7674
rect 7529 7658 7535 7660
rect 7506 7655 7535 7658
rect 7827 7654 7830 7660
rect 7856 7674 7859 7680
rect 8195 7674 8198 7680
rect 7856 7660 8198 7674
rect 7856 7654 7859 7660
rect 8195 7654 8198 7660
rect 8224 7654 8227 7680
rect 8747 7654 8750 7680
rect 8776 7654 8779 7680
rect 19925 7654 19928 7680
rect 19954 7654 19957 7680
rect 21673 7654 21676 7680
rect 21702 7674 21705 7680
rect 22272 7675 22301 7678
rect 22272 7674 22278 7675
rect 21702 7660 22278 7674
rect 21702 7654 21705 7660
rect 22272 7658 22278 7660
rect 22295 7658 22301 7675
rect 22272 7655 22301 7658
rect 22916 7675 22945 7678
rect 22916 7658 22922 7675
rect 22939 7674 22945 7675
rect 24341 7674 24344 7680
rect 22939 7660 24344 7674
rect 22939 7658 22945 7660
rect 22916 7655 22945 7658
rect 24341 7654 24344 7660
rect 24370 7654 24373 7680
rect 26819 7674 26833 7694
rect 26871 7688 26874 7714
rect 26900 7713 26924 7714
rect 26947 7733 26976 7736
rect 26947 7716 26953 7733
rect 26970 7716 26976 7733
rect 26995 7726 27001 7743
rect 27018 7742 27024 7743
rect 27046 7743 27075 7746
rect 27018 7726 27032 7742
rect 26995 7723 27032 7726
rect 27046 7726 27052 7743
rect 27069 7742 27075 7743
rect 27101 7742 27104 7748
rect 27069 7728 27104 7742
rect 27069 7726 27075 7728
rect 27046 7723 27075 7726
rect 26947 7713 26976 7716
rect 26900 7694 26917 7713
rect 26900 7688 26903 7694
rect 26952 7674 26966 7713
rect 27018 7708 27032 7723
rect 27101 7722 27104 7728
rect 27130 7722 27133 7748
rect 27930 7743 27959 7746
rect 27930 7726 27936 7743
rect 27953 7742 27959 7743
rect 27975 7742 27978 7748
rect 27953 7728 27978 7742
rect 27953 7726 27959 7728
rect 27930 7723 27959 7726
rect 27975 7722 27978 7728
rect 28004 7722 28007 7748
rect 28067 7722 28070 7748
rect 28096 7746 28099 7748
rect 28096 7743 28114 7746
rect 28108 7726 28114 7743
rect 28619 7742 28622 7748
rect 28096 7723 28114 7726
rect 28260 7728 28622 7742
rect 28096 7722 28099 7723
rect 27745 7708 27748 7714
rect 27018 7694 27748 7708
rect 27745 7688 27748 7694
rect 27774 7688 27777 7714
rect 27883 7688 27886 7714
rect 27912 7708 27915 7714
rect 28129 7709 28158 7712
rect 28129 7708 28135 7709
rect 27912 7694 28135 7708
rect 27912 7688 27915 7694
rect 28129 7692 28135 7694
rect 28152 7708 28158 7709
rect 28260 7708 28274 7728
rect 28619 7722 28622 7728
rect 28648 7722 28651 7748
rect 29309 7722 29312 7748
rect 29338 7742 29341 7748
rect 29494 7743 29523 7746
rect 29494 7742 29500 7743
rect 29338 7728 29500 7742
rect 29338 7722 29341 7728
rect 29494 7726 29500 7728
rect 29517 7726 29523 7743
rect 29494 7723 29523 7726
rect 29539 7722 29542 7748
rect 29568 7722 29571 7748
rect 29723 7722 29726 7748
rect 29752 7722 29755 7748
rect 28152 7694 28274 7708
rect 28152 7692 28158 7694
rect 28129 7689 28158 7692
rect 29401 7688 29404 7714
rect 29430 7708 29433 7714
rect 29632 7709 29661 7712
rect 29632 7708 29638 7709
rect 29430 7694 29638 7708
rect 29430 7688 29433 7694
rect 29632 7692 29638 7694
rect 29655 7692 29661 7709
rect 29632 7689 29661 7692
rect 29677 7688 29680 7714
rect 29706 7688 29709 7714
rect 27285 7674 27288 7680
rect 26819 7660 27288 7674
rect 27285 7654 27288 7660
rect 27314 7654 27317 7680
rect 3036 7592 29992 7640
rect 6126 7573 6155 7576
rect 6126 7556 6132 7573
rect 6149 7572 6155 7573
rect 6171 7572 6174 7578
rect 6149 7558 6174 7572
rect 6149 7556 6155 7558
rect 6126 7553 6155 7556
rect 6171 7552 6174 7558
rect 6200 7552 6203 7578
rect 15510 7573 15539 7576
rect 15510 7556 15516 7573
rect 15533 7572 15539 7573
rect 15785 7572 15788 7578
rect 15533 7558 15788 7572
rect 15533 7556 15539 7558
rect 15510 7553 15539 7556
rect 15785 7552 15788 7558
rect 15814 7552 15817 7578
rect 18269 7552 18272 7578
rect 18298 7552 18301 7578
rect 21443 7572 21446 7578
rect 20394 7558 21446 7572
rect 5987 7518 5990 7544
rect 6016 7538 6019 7544
rect 6034 7539 6063 7542
rect 6034 7538 6040 7539
rect 6016 7524 6040 7538
rect 6016 7518 6019 7524
rect 6034 7522 6040 7524
rect 6057 7538 6063 7539
rect 6079 7538 6082 7544
rect 6057 7524 6082 7538
rect 6057 7522 6063 7524
rect 6034 7519 6063 7522
rect 6079 7518 6082 7524
rect 6108 7518 6111 7544
rect 7137 7518 7140 7544
rect 7166 7518 7169 7544
rect 7689 7518 7692 7544
rect 7718 7538 7721 7544
rect 8058 7539 8087 7542
rect 8058 7538 8064 7539
rect 7718 7524 8064 7538
rect 7718 7518 7721 7524
rect 8058 7522 8064 7524
rect 8081 7522 8087 7539
rect 8058 7519 8087 7522
rect 9346 7539 9375 7542
rect 9346 7522 9352 7539
rect 9369 7538 9375 7539
rect 9691 7539 9720 7542
rect 9691 7538 9697 7539
rect 9369 7524 9697 7538
rect 9369 7522 9375 7524
rect 9346 7519 9375 7522
rect 9691 7522 9697 7524
rect 9714 7522 9720 7539
rect 11645 7538 11648 7544
rect 9691 7519 9720 7522
rect 10366 7524 10518 7538
rect 6172 7505 6201 7508
rect 6172 7488 6178 7505
rect 6195 7504 6201 7505
rect 6217 7504 6220 7510
rect 6195 7490 6220 7504
rect 6195 7488 6201 7490
rect 6172 7485 6201 7488
rect 6217 7484 6220 7490
rect 6246 7484 6249 7510
rect 7643 7484 7646 7510
rect 7672 7504 7675 7510
rect 7920 7505 7949 7508
rect 7920 7504 7926 7505
rect 7672 7490 7926 7504
rect 7672 7484 7675 7490
rect 7920 7488 7926 7490
rect 7943 7504 7949 7505
rect 9069 7504 9072 7510
rect 7943 7490 9072 7504
rect 7943 7488 7949 7490
rect 7920 7485 7949 7488
rect 9069 7484 9072 7490
rect 9098 7484 9101 7510
rect 9253 7484 9256 7510
rect 9282 7484 9285 7510
rect 9392 7505 9421 7508
rect 9392 7488 9398 7505
rect 9415 7504 9421 7505
rect 9437 7504 9440 7510
rect 9415 7490 9440 7504
rect 9415 7488 9421 7490
rect 9392 7485 9421 7488
rect 9437 7484 9440 7490
rect 9466 7484 9469 7510
rect 9575 7484 9578 7510
rect 9604 7504 9607 7510
rect 9640 7505 9669 7508
rect 9640 7504 9646 7505
rect 9604 7490 9646 7504
rect 9604 7484 9607 7490
rect 9640 7488 9646 7490
rect 9663 7504 9669 7505
rect 10366 7504 10380 7524
rect 9663 7490 10380 7504
rect 9663 7488 9669 7490
rect 9640 7485 9669 7488
rect 10403 7484 10406 7510
rect 10432 7484 10435 7510
rect 10504 7508 10518 7524
rect 10734 7524 11648 7538
rect 10734 7508 10748 7524
rect 11645 7518 11648 7524
rect 11674 7518 11677 7544
rect 19236 7539 19265 7542
rect 19236 7522 19242 7539
rect 19259 7538 19265 7539
rect 19649 7538 19652 7544
rect 19259 7524 19652 7538
rect 19259 7522 19265 7524
rect 19236 7519 19265 7522
rect 19649 7518 19652 7524
rect 19678 7518 19681 7544
rect 10496 7505 10525 7508
rect 10496 7488 10502 7505
rect 10519 7504 10525 7505
rect 10726 7505 10755 7508
rect 10726 7504 10732 7505
rect 10519 7490 10732 7504
rect 10519 7488 10525 7490
rect 10496 7485 10525 7488
rect 10726 7488 10732 7490
rect 10749 7488 10755 7505
rect 10726 7485 10755 7488
rect 10818 7505 10847 7508
rect 10818 7488 10824 7505
rect 10841 7488 10847 7505
rect 10818 7485 10847 7488
rect 10864 7505 10893 7508
rect 10864 7488 10870 7505
rect 10887 7504 10893 7505
rect 11093 7504 11096 7510
rect 10887 7490 11096 7504
rect 10887 7488 10893 7490
rect 10864 7485 10893 7488
rect 10826 7470 10840 7485
rect 11093 7484 11096 7490
rect 11122 7504 11125 7510
rect 11507 7504 11510 7510
rect 11122 7490 11510 7504
rect 11122 7484 11125 7490
rect 11507 7484 11510 7490
rect 11536 7504 11539 7510
rect 11554 7505 11583 7508
rect 11554 7504 11560 7505
rect 11536 7490 11560 7504
rect 11536 7484 11539 7490
rect 11554 7488 11560 7490
rect 11577 7488 11583 7505
rect 11554 7485 11583 7488
rect 11692 7505 11721 7508
rect 11692 7488 11698 7505
rect 11715 7504 11721 7505
rect 11829 7504 11832 7510
rect 11715 7490 11832 7504
rect 11715 7488 11721 7490
rect 11692 7485 11721 7488
rect 11700 7470 11714 7485
rect 11829 7484 11832 7490
rect 11858 7484 11861 7510
rect 15326 7505 15355 7508
rect 15326 7488 15332 7505
rect 15349 7504 15355 7505
rect 15739 7504 15742 7510
rect 15349 7490 15742 7504
rect 15349 7488 15355 7490
rect 15326 7485 15355 7488
rect 15739 7484 15742 7490
rect 15768 7484 15771 7510
rect 18224 7505 18253 7508
rect 18224 7488 18230 7505
rect 18247 7488 18253 7505
rect 18224 7485 18253 7488
rect 10826 7456 11714 7470
rect 14313 7450 14316 7476
rect 14342 7470 14345 7476
rect 15280 7471 15309 7474
rect 15280 7470 15286 7471
rect 14342 7456 15286 7470
rect 14342 7450 14345 7456
rect 15280 7454 15286 7456
rect 15303 7454 15309 7471
rect 18232 7470 18246 7485
rect 18315 7484 18318 7510
rect 18344 7484 18347 7510
rect 18959 7484 18962 7510
rect 18988 7484 18991 7510
rect 19097 7484 19100 7510
rect 19126 7484 19129 7510
rect 19327 7484 19330 7510
rect 19356 7504 19359 7510
rect 20110 7505 20139 7508
rect 20110 7504 20116 7505
rect 19356 7490 20116 7504
rect 19356 7484 19359 7490
rect 20110 7488 20116 7490
rect 20133 7488 20139 7505
rect 20110 7485 20139 7488
rect 20339 7484 20342 7510
rect 20368 7504 20371 7510
rect 20394 7508 20408 7558
rect 21443 7552 21446 7558
rect 21472 7552 21475 7578
rect 24319 7573 24348 7576
rect 24319 7556 24325 7573
rect 24342 7572 24348 7573
rect 24479 7572 24482 7578
rect 24342 7558 24482 7572
rect 24342 7556 24348 7558
rect 24319 7553 24348 7556
rect 24479 7552 24482 7558
rect 24508 7552 24511 7578
rect 26871 7576 26874 7578
rect 26849 7573 26874 7576
rect 26849 7556 26855 7573
rect 26872 7556 26874 7573
rect 26849 7553 26874 7556
rect 26871 7552 26874 7553
rect 26900 7552 26903 7578
rect 29149 7573 29178 7576
rect 29149 7556 29155 7573
rect 29172 7572 29178 7573
rect 29539 7572 29542 7578
rect 29172 7558 29542 7572
rect 29172 7556 29178 7558
rect 29149 7553 29178 7556
rect 29539 7552 29542 7558
rect 29568 7552 29571 7578
rect 20478 7539 20507 7542
rect 20478 7522 20484 7539
rect 20501 7538 20507 7539
rect 20501 7524 20707 7538
rect 20501 7522 20507 7524
rect 20478 7519 20507 7522
rect 20386 7505 20415 7508
rect 20386 7504 20392 7505
rect 20368 7490 20392 7504
rect 20368 7484 20371 7490
rect 20386 7488 20392 7490
rect 20409 7488 20415 7505
rect 20386 7485 20415 7488
rect 18968 7470 18982 7484
rect 18232 7456 18982 7470
rect 15280 7451 15309 7454
rect 7966 7437 7995 7440
rect 7966 7420 7972 7437
rect 7989 7436 7995 7437
rect 8195 7436 8198 7442
rect 7989 7422 8198 7436
rect 7989 7420 7995 7422
rect 7966 7417 7995 7420
rect 8195 7416 8198 7422
rect 8224 7416 8227 7442
rect 9115 7416 9118 7442
rect 9144 7436 9147 7442
rect 9254 7437 9283 7440
rect 9254 7436 9260 7437
rect 9144 7422 9260 7436
rect 9144 7416 9147 7422
rect 9254 7420 9260 7422
rect 9277 7420 9283 7437
rect 9254 7417 9283 7420
rect 10587 7416 10590 7442
rect 10616 7436 10619 7442
rect 10616 7422 10978 7436
rect 10616 7416 10619 7422
rect 6034 7403 6063 7406
rect 6034 7386 6040 7403
rect 6057 7402 6063 7403
rect 6125 7402 6128 7408
rect 6057 7388 6128 7402
rect 6057 7386 6063 7388
rect 6034 7383 6063 7386
rect 6125 7382 6128 7388
rect 6154 7382 6157 7408
rect 6585 7382 6588 7408
rect 6614 7402 6617 7408
rect 6861 7402 6864 7408
rect 6614 7388 6864 7402
rect 6614 7382 6617 7388
rect 6861 7382 6864 7388
rect 6890 7402 6893 7408
rect 7184 7403 7213 7406
rect 7184 7402 7190 7403
rect 6890 7388 7190 7402
rect 6890 7382 6893 7388
rect 7184 7386 7190 7388
rect 7207 7402 7213 7403
rect 7597 7402 7600 7408
rect 7207 7388 7600 7402
rect 7207 7386 7213 7388
rect 7184 7383 7213 7386
rect 7597 7382 7600 7388
rect 7626 7382 7629 7408
rect 7735 7382 7738 7408
rect 7764 7402 7767 7408
rect 7920 7403 7949 7406
rect 7920 7402 7926 7403
rect 7764 7388 7926 7402
rect 7764 7382 7767 7388
rect 7920 7386 7926 7388
rect 7943 7386 7949 7403
rect 7920 7383 7949 7386
rect 10403 7382 10406 7408
rect 10432 7382 10435 7408
rect 10725 7382 10728 7408
rect 10754 7382 10757 7408
rect 10964 7406 10978 7422
rect 11553 7416 11556 7442
rect 11582 7416 11585 7442
rect 20693 7436 20707 7524
rect 20753 7518 20756 7544
rect 20782 7518 20785 7544
rect 21029 7518 21032 7544
rect 21058 7518 21061 7544
rect 21075 7518 21078 7544
rect 21104 7518 21107 7544
rect 23513 7542 23516 7544
rect 23491 7539 23516 7542
rect 23491 7538 23497 7539
rect 22740 7524 23497 7538
rect 20983 7484 20986 7510
rect 21012 7484 21015 7510
rect 20800 7471 20829 7474
rect 20800 7454 20806 7471
rect 20823 7470 20829 7471
rect 22685 7470 22688 7476
rect 20823 7456 22688 7470
rect 20823 7454 20829 7456
rect 20800 7451 20829 7454
rect 22685 7450 22688 7456
rect 22714 7450 22717 7476
rect 21397 7436 21400 7442
rect 20693 7422 21400 7436
rect 21397 7416 21400 7422
rect 21426 7416 21429 7442
rect 10956 7403 10985 7406
rect 10956 7386 10962 7403
rect 10979 7386 10985 7403
rect 10956 7383 10985 7386
rect 20707 7382 20710 7408
rect 20736 7402 20739 7408
rect 22740 7402 22754 7524
rect 23491 7522 23497 7524
rect 23514 7522 23516 7539
rect 23491 7519 23516 7522
rect 23513 7518 23516 7519
rect 23542 7518 23545 7544
rect 25859 7518 25862 7544
rect 25888 7538 25891 7544
rect 26025 7539 26054 7542
rect 26025 7538 26031 7539
rect 25888 7524 26031 7538
rect 25888 7518 25891 7524
rect 26025 7522 26031 7524
rect 26048 7538 26054 7539
rect 26089 7538 26092 7544
rect 26048 7524 26092 7538
rect 26048 7522 26054 7524
rect 26025 7519 26054 7522
rect 26089 7518 26092 7524
rect 26118 7518 26121 7544
rect 28343 7542 28346 7544
rect 28325 7539 28346 7542
rect 28325 7522 28331 7539
rect 28325 7519 28346 7522
rect 28343 7518 28346 7519
rect 28372 7518 28375 7544
rect 23237 7484 23240 7510
rect 23266 7504 23269 7510
rect 23284 7505 23313 7508
rect 23284 7504 23290 7505
rect 23266 7490 23290 7504
rect 23266 7484 23269 7490
rect 23284 7488 23290 7490
rect 23307 7488 23313 7505
rect 23284 7485 23313 7488
rect 23445 7505 23474 7508
rect 23445 7488 23451 7505
rect 23468 7504 23474 7505
rect 23559 7504 23562 7510
rect 23468 7490 23562 7504
rect 23468 7488 23474 7490
rect 23445 7485 23474 7488
rect 23559 7484 23562 7490
rect 23588 7484 23591 7510
rect 25975 7505 26004 7508
rect 25975 7488 25981 7505
rect 25998 7504 26004 7505
rect 26135 7504 26138 7510
rect 25998 7490 26138 7504
rect 25998 7488 26004 7490
rect 25975 7485 26004 7488
rect 26135 7484 26138 7490
rect 26164 7484 26167 7510
rect 27975 7484 27978 7510
rect 28004 7504 28007 7510
rect 28114 7505 28143 7508
rect 28114 7504 28120 7505
rect 28004 7490 28120 7504
rect 28004 7484 28007 7490
rect 28114 7488 28120 7490
rect 28137 7488 28143 7505
rect 28114 7485 28143 7488
rect 28275 7505 28304 7508
rect 28275 7488 28281 7505
rect 28298 7504 28304 7505
rect 28389 7504 28392 7510
rect 28298 7490 28392 7504
rect 28298 7488 28304 7490
rect 28275 7485 28304 7488
rect 28389 7484 28392 7490
rect 28418 7484 28421 7510
rect 25813 7450 25816 7476
rect 25842 7450 25845 7476
rect 20736 7388 22754 7402
rect 20736 7382 20739 7388
rect 23513 7382 23516 7408
rect 23542 7402 23545 7408
rect 24663 7402 24666 7408
rect 23542 7388 24666 7402
rect 23542 7382 23545 7388
rect 24663 7382 24666 7388
rect 24692 7382 24695 7408
rect 3036 7320 29992 7368
rect 8793 7280 8796 7306
rect 8822 7300 8825 7306
rect 8840 7301 8869 7304
rect 8840 7300 8846 7301
rect 8822 7286 8846 7300
rect 8822 7280 8825 7286
rect 8840 7284 8846 7286
rect 8863 7284 8869 7301
rect 8840 7281 8869 7284
rect 9069 7280 9072 7306
rect 9098 7280 9101 7306
rect 10403 7280 10406 7306
rect 10432 7300 10435 7306
rect 10763 7301 10792 7304
rect 10763 7300 10769 7301
rect 10432 7286 10769 7300
rect 10432 7280 10435 7286
rect 10763 7284 10769 7286
rect 10786 7284 10792 7301
rect 10763 7281 10792 7284
rect 14313 7280 14316 7306
rect 14342 7280 14345 7306
rect 21075 7280 21078 7306
rect 21104 7300 21107 7306
rect 23237 7300 23240 7306
rect 21104 7286 23240 7300
rect 21104 7280 21107 7286
rect 23237 7280 23240 7286
rect 23266 7280 23269 7306
rect 25675 7280 25678 7306
rect 25704 7300 25707 7306
rect 25813 7300 25816 7306
rect 25704 7286 25816 7300
rect 25704 7280 25707 7286
rect 25813 7280 25816 7286
rect 25842 7300 25845 7306
rect 25842 7286 27676 7300
rect 25842 7280 25845 7286
rect 10587 7266 10590 7272
rect 8986 7252 10590 7266
rect 6171 7212 6174 7238
rect 6200 7232 6203 7238
rect 6540 7233 6569 7236
rect 6540 7232 6546 7233
rect 6200 7218 6546 7232
rect 6200 7212 6203 7218
rect 6540 7216 6546 7218
rect 6563 7216 6569 7233
rect 6540 7213 6569 7216
rect 7597 7212 7600 7238
rect 7626 7212 7629 7238
rect 7735 7212 7738 7238
rect 7764 7212 7767 7238
rect 8103 7212 8106 7238
rect 8132 7232 8135 7238
rect 8610 7233 8639 7236
rect 8610 7232 8616 7233
rect 8132 7218 8616 7232
rect 8132 7212 8135 7218
rect 8610 7216 8616 7218
rect 8633 7232 8639 7233
rect 8633 7218 8954 7232
rect 8633 7216 8639 7218
rect 8610 7213 8639 7216
rect 5527 7178 5530 7204
rect 5556 7178 5559 7204
rect 8940 7202 8954 7218
rect 8986 7202 9000 7252
rect 10587 7246 10590 7252
rect 10616 7246 10619 7272
rect 11829 7246 11832 7272
rect 11858 7266 11861 7272
rect 12060 7267 12089 7270
rect 12060 7266 12066 7267
rect 11858 7252 12066 7266
rect 11858 7246 11861 7252
rect 12060 7250 12066 7252
rect 12083 7250 12089 7267
rect 21397 7266 21400 7272
rect 12060 7247 12089 7250
rect 19106 7252 21400 7266
rect 9023 7212 9026 7238
rect 9052 7232 9055 7238
rect 9714 7233 9743 7236
rect 9714 7232 9720 7233
rect 9052 7218 9720 7232
rect 9052 7212 9055 7218
rect 9714 7216 9720 7218
rect 9737 7216 9743 7233
rect 9714 7213 9743 7216
rect 10357 7212 10360 7238
rect 10386 7232 10389 7238
rect 10634 7233 10663 7236
rect 10634 7232 10640 7233
rect 10386 7218 10640 7232
rect 10386 7212 10389 7218
rect 10634 7216 10640 7218
rect 10657 7232 10663 7233
rect 10817 7232 10820 7238
rect 10657 7218 10820 7232
rect 10657 7216 10663 7218
rect 10634 7213 10663 7216
rect 10817 7212 10820 7218
rect 10846 7212 10849 7238
rect 11645 7212 11648 7238
rect 11674 7232 11677 7238
rect 12106 7233 12135 7236
rect 12106 7232 12112 7233
rect 11674 7218 12112 7232
rect 11674 7212 11677 7218
rect 12106 7216 12112 7218
rect 12129 7216 12135 7233
rect 12106 7213 12135 7216
rect 14037 7212 14040 7238
rect 14066 7232 14069 7238
rect 14084 7233 14113 7236
rect 14084 7232 14090 7233
rect 14066 7218 14090 7232
rect 14066 7212 14069 7218
rect 14084 7216 14090 7218
rect 14107 7216 14113 7233
rect 18959 7232 18962 7238
rect 14084 7213 14113 7216
rect 18692 7218 18962 7232
rect 8932 7199 8961 7202
rect 8932 7182 8938 7199
rect 8955 7182 8961 7199
rect 8932 7179 8961 7182
rect 8978 7199 9007 7202
rect 8978 7182 8984 7199
rect 9001 7182 9007 7199
rect 8978 7179 9007 7182
rect 5665 7144 5668 7170
rect 5694 7144 5697 7170
rect 5941 7144 5944 7170
rect 5970 7144 5973 7170
rect 6033 7144 6036 7170
rect 6062 7144 6065 7170
rect 7597 7144 7600 7170
rect 7626 7164 7629 7170
rect 7689 7164 7692 7170
rect 7626 7150 7692 7164
rect 7626 7144 7629 7150
rect 7689 7144 7692 7150
rect 7718 7164 7721 7170
rect 7718 7150 7981 7164
rect 7718 7144 7721 7150
rect 8885 7144 8888 7170
rect 8914 7164 8917 7170
rect 8986 7164 9000 7179
rect 9575 7178 9578 7204
rect 9604 7178 9607 7204
rect 9622 7199 9651 7202
rect 9622 7182 9628 7199
rect 9645 7182 9651 7199
rect 9622 7179 9651 7182
rect 8914 7150 9000 7164
rect 8914 7144 8917 7150
rect 9437 7144 9440 7170
rect 9466 7164 9469 7170
rect 9630 7164 9644 7179
rect 11507 7178 11510 7204
rect 11536 7198 11539 7204
rect 11968 7199 11997 7202
rect 11968 7198 11974 7199
rect 11536 7184 11974 7198
rect 11536 7178 11539 7184
rect 11968 7182 11974 7184
rect 11991 7182 11997 7199
rect 11968 7179 11997 7182
rect 14130 7199 14159 7202
rect 14130 7182 14136 7199
rect 14153 7198 14159 7199
rect 14405 7198 14408 7204
rect 14153 7184 14408 7198
rect 14153 7182 14159 7184
rect 14130 7179 14159 7182
rect 14405 7178 14408 7184
rect 14434 7178 14437 7204
rect 15785 7178 15788 7204
rect 15814 7198 15817 7204
rect 18637 7198 18640 7204
rect 15814 7184 18640 7198
rect 15814 7178 15817 7184
rect 18637 7178 18640 7184
rect 18666 7178 18669 7204
rect 18692 7202 18706 7218
rect 18959 7212 18962 7218
rect 18988 7212 18991 7238
rect 18684 7199 18713 7202
rect 18684 7182 18690 7199
rect 18707 7182 18713 7199
rect 18684 7179 18713 7182
rect 18822 7199 18851 7202
rect 18822 7182 18828 7199
rect 18845 7182 18851 7199
rect 18822 7179 18851 7182
rect 18914 7199 18943 7202
rect 18914 7182 18920 7199
rect 18937 7198 18943 7199
rect 19106 7198 19120 7252
rect 21397 7246 21400 7252
rect 21426 7246 21429 7272
rect 19143 7212 19146 7238
rect 19172 7232 19175 7238
rect 19742 7233 19771 7236
rect 19742 7232 19748 7233
rect 19172 7218 19748 7232
rect 19172 7212 19175 7218
rect 19742 7216 19748 7218
rect 19765 7216 19771 7233
rect 19742 7213 19771 7216
rect 19834 7233 19863 7236
rect 19834 7216 19840 7233
rect 19857 7232 19863 7233
rect 20063 7232 20066 7238
rect 19857 7218 20066 7232
rect 19857 7216 19863 7218
rect 19834 7213 19863 7216
rect 20063 7212 20066 7218
rect 20092 7212 20095 7238
rect 22179 7212 22182 7238
rect 22208 7232 22211 7238
rect 26742 7236 26756 7286
rect 27662 7266 27676 7286
rect 27745 7280 27748 7306
rect 27774 7304 27777 7306
rect 27774 7301 27798 7304
rect 27774 7284 27775 7301
rect 27792 7284 27798 7301
rect 27774 7281 27798 7284
rect 27774 7280 27777 7281
rect 27975 7266 27978 7272
rect 27662 7252 27978 7266
rect 27975 7246 27978 7252
rect 28004 7246 28007 7272
rect 26734 7233 26763 7236
rect 22208 7218 22478 7232
rect 22208 7212 22211 7218
rect 18937 7184 19120 7198
rect 19558 7199 19587 7202
rect 18937 7182 18943 7184
rect 18914 7179 18943 7182
rect 19558 7182 19564 7199
rect 19581 7198 19587 7199
rect 19603 7198 19606 7204
rect 19581 7184 19606 7198
rect 19581 7182 19587 7184
rect 19558 7179 19587 7182
rect 9466 7150 9644 7164
rect 9466 7144 9469 7150
rect 11001 7144 11004 7170
rect 11030 7144 11033 7170
rect 18315 7144 18318 7170
rect 18344 7164 18347 7170
rect 18830 7164 18844 7179
rect 19603 7178 19606 7184
rect 19632 7178 19635 7204
rect 19696 7199 19725 7202
rect 19696 7182 19702 7199
rect 19719 7198 19725 7199
rect 19787 7198 19790 7204
rect 19719 7184 19790 7198
rect 19719 7182 19725 7184
rect 19696 7179 19725 7182
rect 19787 7178 19790 7184
rect 19816 7198 19819 7204
rect 19971 7198 19974 7204
rect 19816 7184 19974 7198
rect 19816 7178 19819 7184
rect 19971 7178 19974 7184
rect 20000 7178 20003 7204
rect 22133 7178 22136 7204
rect 22162 7198 22165 7204
rect 22464 7202 22478 7218
rect 26734 7216 26740 7233
rect 26757 7216 26763 7233
rect 26734 7213 26763 7216
rect 22226 7199 22255 7202
rect 22226 7198 22232 7199
rect 22162 7184 22232 7198
rect 22162 7178 22165 7184
rect 22226 7182 22232 7184
rect 22249 7182 22255 7199
rect 22226 7179 22255 7182
rect 22456 7199 22485 7202
rect 22456 7182 22462 7199
rect 22479 7182 22485 7199
rect 22456 7179 22485 7182
rect 22639 7178 22642 7204
rect 22668 7178 22671 7204
rect 22777 7178 22780 7204
rect 22806 7198 22809 7204
rect 22824 7199 22853 7202
rect 22824 7198 22830 7199
rect 22806 7184 22830 7198
rect 22806 7178 22809 7184
rect 22824 7182 22830 7184
rect 22847 7182 22853 7199
rect 22824 7179 22853 7182
rect 26135 7178 26138 7204
rect 26164 7198 26167 7204
rect 26889 7199 26918 7202
rect 26889 7198 26895 7199
rect 26164 7184 26895 7198
rect 26164 7178 26167 7184
rect 26889 7182 26895 7184
rect 26912 7182 26918 7199
rect 26889 7179 26918 7182
rect 20339 7164 20342 7170
rect 18344 7150 20342 7164
rect 18344 7144 18347 7150
rect 20339 7144 20342 7150
rect 20368 7144 20371 7170
rect 21305 7164 21308 7170
rect 20670 7150 21308 7164
rect 9299 7110 9302 7136
rect 9328 7130 9331 7136
rect 9714 7131 9743 7134
rect 9714 7130 9720 7131
rect 9328 7116 9720 7130
rect 9328 7110 9331 7116
rect 9714 7114 9720 7116
rect 9737 7114 9743 7131
rect 9714 7111 9743 7114
rect 11139 7110 11142 7136
rect 11168 7130 11171 7136
rect 11876 7131 11905 7134
rect 11876 7130 11882 7131
rect 11168 7116 11882 7130
rect 11168 7110 11171 7116
rect 11876 7114 11882 7116
rect 11899 7114 11905 7131
rect 11876 7111 11905 7114
rect 18407 7110 18410 7136
rect 18436 7130 18439 7136
rect 18592 7131 18621 7134
rect 18592 7130 18598 7131
rect 18436 7116 18598 7130
rect 18436 7110 18439 7116
rect 18592 7114 18598 7116
rect 18615 7114 18621 7131
rect 18592 7111 18621 7114
rect 19373 7110 19376 7136
rect 19402 7130 19405 7136
rect 20670 7130 20684 7150
rect 21305 7144 21308 7150
rect 21334 7164 21337 7170
rect 24203 7164 24206 7170
rect 21334 7150 24206 7164
rect 21334 7144 21337 7150
rect 24203 7144 24206 7150
rect 24232 7144 24235 7170
rect 26963 7168 26966 7170
rect 26945 7165 26966 7168
rect 26945 7148 26951 7165
rect 26945 7145 26966 7148
rect 26963 7144 26966 7145
rect 26992 7144 26995 7170
rect 19402 7116 20684 7130
rect 19402 7110 19405 7116
rect 21121 7110 21124 7136
rect 21150 7130 21153 7136
rect 21213 7130 21216 7136
rect 21150 7116 21216 7130
rect 21150 7110 21153 7116
rect 21213 7110 21216 7116
rect 21242 7130 21245 7136
rect 21443 7130 21446 7136
rect 21242 7116 21446 7130
rect 21242 7110 21245 7116
rect 21443 7110 21446 7116
rect 21472 7110 21475 7136
rect 22364 7131 22393 7134
rect 22364 7114 22370 7131
rect 22387 7130 22393 7131
rect 22593 7130 22596 7136
rect 22387 7116 22596 7130
rect 22387 7114 22393 7116
rect 22364 7111 22393 7114
rect 22593 7110 22596 7116
rect 22622 7110 22625 7136
rect 22915 7110 22918 7136
rect 22944 7130 22947 7136
rect 24893 7130 24896 7136
rect 22944 7116 24896 7130
rect 22944 7110 22947 7116
rect 24893 7110 24896 7116
rect 24922 7110 24925 7136
rect 3036 7048 29992 7096
rect 5665 7008 5668 7034
rect 5694 7028 5697 7034
rect 6034 7029 6063 7032
rect 6034 7028 6040 7029
rect 5694 7014 6040 7028
rect 5694 7008 5697 7014
rect 6034 7012 6040 7014
rect 6057 7012 6063 7029
rect 6034 7009 6063 7012
rect 8288 7029 8317 7032
rect 8288 7012 8294 7029
rect 8311 7028 8317 7029
rect 8793 7028 8796 7034
rect 8311 7014 8796 7028
rect 8311 7012 8317 7014
rect 8288 7009 8317 7012
rect 8793 7008 8796 7014
rect 8822 7008 8825 7034
rect 10725 7008 10728 7034
rect 10754 7028 10757 7034
rect 11048 7029 11077 7032
rect 11048 7028 11054 7029
rect 10754 7014 11054 7028
rect 10754 7008 10757 7014
rect 11048 7012 11054 7014
rect 11071 7012 11077 7029
rect 14452 7029 14481 7032
rect 14452 7028 14458 7029
rect 11048 7009 11077 7012
rect 13724 7014 14458 7028
rect 10449 6974 10452 7000
rect 10478 6994 10481 7000
rect 13724 6998 13738 7014
rect 14452 7012 14458 7014
rect 14475 7012 14481 7029
rect 14452 7009 14481 7012
rect 20386 7029 20415 7032
rect 20386 7012 20392 7029
rect 20409 7028 20415 7029
rect 21121 7028 21124 7034
rect 20409 7014 21124 7028
rect 20409 7012 20415 7014
rect 20386 7009 20415 7012
rect 21121 7008 21124 7014
rect 21150 7008 21153 7034
rect 22111 7029 22140 7032
rect 22111 7012 22117 7029
rect 22134 7028 22140 7029
rect 22134 7014 22877 7028
rect 22134 7012 22140 7014
rect 22111 7009 22140 7012
rect 10956 6995 10985 6998
rect 10956 6994 10962 6995
rect 10478 6980 10962 6994
rect 10478 6974 10481 6980
rect 10956 6978 10962 6980
rect 10979 6978 10985 6995
rect 10956 6975 10985 6978
rect 13716 6995 13745 6998
rect 13716 6978 13722 6995
rect 13739 6978 13745 6995
rect 13716 6975 13745 6978
rect 13807 6974 13810 7000
rect 13836 6994 13839 7000
rect 13836 6980 14382 6994
rect 13836 6974 13839 6980
rect 6125 6940 6128 6966
rect 6154 6940 6157 6966
rect 8103 6940 8106 6966
rect 8132 6960 8135 6966
rect 8196 6961 8225 6964
rect 8196 6960 8202 6961
rect 8132 6946 8202 6960
rect 8132 6940 8135 6946
rect 8196 6944 8202 6946
rect 8219 6944 8225 6961
rect 8196 6941 8225 6944
rect 8334 6961 8363 6964
rect 8334 6944 8340 6961
rect 8357 6960 8363 6961
rect 8885 6960 8888 6966
rect 8357 6946 8888 6960
rect 8357 6944 8363 6946
rect 8334 6941 8363 6944
rect 8885 6940 8888 6946
rect 8914 6940 8917 6966
rect 11094 6961 11123 6964
rect 11094 6944 11100 6961
rect 11117 6960 11123 6961
rect 11829 6960 11832 6966
rect 11117 6946 11832 6960
rect 11117 6944 11123 6946
rect 11094 6941 11123 6944
rect 11829 6940 11832 6946
rect 11858 6940 11861 6966
rect 13854 6961 13883 6964
rect 13854 6944 13860 6961
rect 13877 6960 13883 6961
rect 14267 6960 14270 6966
rect 13877 6946 14270 6960
rect 13877 6944 13883 6946
rect 13854 6941 13883 6944
rect 14267 6940 14270 6946
rect 14296 6940 14299 6966
rect 14368 6964 14382 6980
rect 15739 6974 15742 7000
rect 15768 6994 15771 7000
rect 18407 6994 18410 7000
rect 15768 6980 18410 6994
rect 15768 6974 15771 6980
rect 14360 6961 14389 6964
rect 14360 6944 14366 6961
rect 14383 6944 14389 6961
rect 15785 6960 15788 6966
rect 14360 6941 14389 6944
rect 14414 6946 15788 6960
rect 6264 6927 6293 6930
rect 6264 6926 6270 6927
rect 6134 6912 6270 6926
rect 6134 6898 6148 6912
rect 6264 6910 6270 6912
rect 6287 6910 6293 6927
rect 6264 6907 6293 6910
rect 14314 6927 14343 6930
rect 14314 6910 14320 6927
rect 14337 6910 14343 6927
rect 14314 6907 14343 6910
rect 6125 6872 6128 6898
rect 6154 6872 6157 6898
rect 8195 6872 8198 6898
rect 8224 6872 8227 6898
rect 10956 6893 10985 6896
rect 10956 6876 10962 6893
rect 10979 6892 10985 6893
rect 11507 6892 11510 6898
rect 10979 6878 11510 6892
rect 10979 6876 10985 6878
rect 10956 6873 10985 6876
rect 11507 6872 11510 6878
rect 11536 6872 11539 6898
rect 14322 6892 14336 6907
rect 14414 6898 14428 6946
rect 15785 6940 15788 6946
rect 15814 6940 15817 6966
rect 16291 6940 16294 6966
rect 16320 6940 16323 6966
rect 17855 6940 17858 6966
rect 17884 6960 17887 6966
rect 18002 6964 18016 6980
rect 18407 6974 18410 6980
rect 18436 6974 18439 7000
rect 20155 6974 20158 7000
rect 20184 6994 20187 7000
rect 21305 6998 21308 7000
rect 21287 6995 21308 6998
rect 20184 6980 21190 6994
rect 20184 6974 20187 6980
rect 17948 6961 17977 6964
rect 17948 6960 17954 6961
rect 17884 6946 17954 6960
rect 17884 6940 17887 6946
rect 17948 6944 17954 6946
rect 17971 6944 17977 6961
rect 17948 6941 17977 6944
rect 17994 6961 18023 6964
rect 17994 6944 18000 6961
rect 18017 6944 18023 6961
rect 17994 6941 18023 6944
rect 18085 6940 18088 6966
rect 18114 6940 18117 6966
rect 18315 6940 18318 6966
rect 18344 6940 18347 6966
rect 19603 6940 19606 6966
rect 19632 6960 19635 6966
rect 19879 6960 19882 6966
rect 19632 6946 19882 6960
rect 19632 6940 19635 6946
rect 19879 6940 19882 6946
rect 19908 6960 19911 6966
rect 20110 6961 20139 6964
rect 20110 6960 20116 6961
rect 19908 6946 20116 6960
rect 19908 6940 19911 6946
rect 20110 6944 20116 6946
rect 20133 6944 20139 6961
rect 20110 6941 20139 6944
rect 20248 6961 20277 6964
rect 20248 6944 20254 6961
rect 20271 6944 20277 6961
rect 20248 6941 20277 6944
rect 14452 6927 14481 6930
rect 14452 6910 14458 6927
rect 14475 6926 14481 6927
rect 14475 6912 15164 6926
rect 14475 6910 14481 6912
rect 14452 6907 14481 6910
rect 14405 6892 14408 6898
rect 14322 6878 14408 6892
rect 14405 6872 14408 6878
rect 14434 6872 14437 6898
rect 15150 6892 15164 6912
rect 15739 6906 15742 6932
rect 15768 6906 15771 6932
rect 15970 6927 15999 6930
rect 15970 6910 15976 6927
rect 15993 6926 15999 6927
rect 16246 6927 16275 6930
rect 16246 6926 16252 6927
rect 15993 6912 16252 6926
rect 15993 6910 15999 6912
rect 15970 6907 15999 6910
rect 16246 6910 16252 6912
rect 16269 6910 16275 6927
rect 16567 6926 16570 6932
rect 16246 6907 16275 6910
rect 16438 6912 16570 6926
rect 16438 6892 16452 6912
rect 16567 6906 16570 6912
rect 16596 6906 16599 6932
rect 18867 6906 18870 6932
rect 18896 6926 18899 6932
rect 19373 6926 19376 6932
rect 18896 6912 19376 6926
rect 18896 6906 18899 6912
rect 19373 6906 19376 6912
rect 19402 6906 19405 6932
rect 19971 6906 19974 6932
rect 20000 6926 20003 6932
rect 20256 6926 20270 6941
rect 20339 6940 20342 6966
rect 20368 6940 20371 6966
rect 21075 6940 21078 6966
rect 21104 6940 21107 6966
rect 21176 6960 21190 6980
rect 21287 6978 21293 6995
rect 21287 6975 21308 6978
rect 21305 6974 21308 6975
rect 21334 6974 21337 7000
rect 22863 6975 22877 7014
rect 23513 6998 23516 7000
rect 23495 6995 23516 6998
rect 23495 6978 23501 6995
rect 23495 6975 23516 6978
rect 22855 6972 22884 6975
rect 23513 6974 23516 6975
rect 23542 6974 23545 7000
rect 25887 6995 25916 6998
rect 25887 6978 25893 6995
rect 25910 6994 25916 6995
rect 25951 6994 25954 7000
rect 25910 6980 25954 6994
rect 25910 6978 25916 6980
rect 25887 6975 25916 6978
rect 25951 6974 25954 6980
rect 25980 6974 25983 7000
rect 29125 6974 29128 7000
rect 29154 6974 29157 7000
rect 21231 6961 21260 6964
rect 21231 6960 21237 6961
rect 21176 6946 21237 6960
rect 21231 6944 21237 6946
rect 21254 6960 21260 6961
rect 21351 6960 21354 6966
rect 21254 6946 21354 6960
rect 21254 6944 21260 6946
rect 21231 6941 21260 6944
rect 21351 6940 21354 6946
rect 21380 6940 21383 6966
rect 22593 6940 22596 6966
rect 22622 6940 22625 6966
rect 22639 6940 22642 6966
rect 22668 6964 22671 6966
rect 22668 6961 22680 6964
rect 22674 6944 22680 6961
rect 22668 6941 22680 6944
rect 22668 6940 22671 6941
rect 22731 6940 22734 6966
rect 22760 6964 22763 6966
rect 22760 6961 22781 6964
rect 22775 6944 22781 6961
rect 22760 6941 22781 6944
rect 22800 6961 22829 6964
rect 22800 6944 22806 6961
rect 22823 6944 22829 6961
rect 22855 6955 22861 6972
rect 22878 6955 22884 6972
rect 22915 6964 22918 6966
rect 22855 6952 22884 6955
rect 22906 6961 22918 6964
rect 22800 6941 22829 6944
rect 22906 6944 22912 6961
rect 22906 6941 22918 6944
rect 22760 6940 22763 6941
rect 20000 6912 20270 6926
rect 20000 6906 20003 6912
rect 22801 6898 22815 6941
rect 22915 6940 22918 6941
rect 22944 6940 22947 6966
rect 23237 6940 23240 6966
rect 23266 6960 23269 6966
rect 23284 6961 23313 6964
rect 23284 6960 23290 6961
rect 23266 6946 23290 6960
rect 23266 6940 23269 6946
rect 23284 6944 23290 6946
rect 23307 6944 23313 6961
rect 23284 6941 23313 6944
rect 23445 6961 23474 6964
rect 23445 6944 23451 6961
rect 23468 6960 23474 6961
rect 23559 6960 23562 6966
rect 23468 6946 23562 6960
rect 23468 6944 23474 6946
rect 23445 6941 23474 6944
rect 23559 6940 23562 6946
rect 23588 6960 23591 6966
rect 23588 6946 24157 6960
rect 23588 6940 23591 6946
rect 24143 6926 24157 6946
rect 24755 6940 24758 6966
rect 24784 6940 24787 6966
rect 24847 6940 24850 6966
rect 24876 6940 24879 6966
rect 24893 6940 24896 6966
rect 24922 6940 24925 6966
rect 25837 6961 25866 6964
rect 25837 6960 25843 6961
rect 24948 6946 25843 6960
rect 24948 6926 24962 6946
rect 25837 6944 25843 6946
rect 25860 6960 25866 6961
rect 26089 6960 26092 6966
rect 25860 6946 26092 6960
rect 25860 6944 25866 6946
rect 25837 6941 25866 6944
rect 26089 6940 26092 6946
rect 26118 6940 26121 6966
rect 29033 6940 29036 6966
rect 29062 6940 29065 6966
rect 29171 6940 29174 6966
rect 29200 6940 29203 6966
rect 29218 6961 29247 6964
rect 29218 6944 29224 6961
rect 29241 6960 29247 6961
rect 29355 6960 29358 6966
rect 29241 6946 29358 6960
rect 29241 6944 29247 6946
rect 29218 6941 29247 6944
rect 29355 6940 29358 6946
rect 29384 6940 29387 6966
rect 24143 6912 24962 6926
rect 15150 6878 16452 6892
rect 16476 6893 16505 6896
rect 16476 6876 16482 6893
rect 16499 6892 16505 6893
rect 17395 6892 17398 6898
rect 16499 6878 17398 6892
rect 16499 6876 16505 6878
rect 16476 6873 16505 6876
rect 17395 6872 17398 6878
rect 17424 6872 17427 6898
rect 22087 6872 22090 6898
rect 22116 6892 22119 6898
rect 22594 6893 22623 6896
rect 22594 6892 22600 6893
rect 22116 6878 22600 6892
rect 22116 6872 22119 6878
rect 22594 6876 22600 6878
rect 22617 6876 22623 6893
rect 22594 6873 22623 6876
rect 22777 6872 22780 6898
rect 22806 6878 22815 6898
rect 22806 6872 22809 6878
rect 6217 6838 6220 6864
rect 6246 6858 6249 6864
rect 6769 6858 6772 6864
rect 6246 6844 6772 6858
rect 6246 6838 6249 6844
rect 6769 6838 6772 6844
rect 6798 6838 6801 6864
rect 13716 6859 13745 6862
rect 13716 6842 13722 6859
rect 13739 6858 13745 6859
rect 13761 6858 13764 6864
rect 13739 6844 13764 6858
rect 13739 6842 13745 6844
rect 13716 6839 13745 6842
rect 13761 6838 13764 6844
rect 13790 6838 13793 6864
rect 24111 6838 24114 6864
rect 24140 6858 24143 6864
rect 24166 6858 24180 6912
rect 25675 6906 25678 6932
rect 25704 6906 25707 6932
rect 24709 6872 24712 6898
rect 24738 6892 24741 6898
rect 26733 6896 26736 6898
rect 24756 6893 24785 6896
rect 24756 6892 24762 6893
rect 24738 6878 24762 6892
rect 24738 6872 24741 6878
rect 24756 6876 24762 6878
rect 24779 6876 24785 6893
rect 24756 6873 24785 6876
rect 26711 6893 26736 6896
rect 26711 6876 26717 6893
rect 26734 6876 26736 6893
rect 26711 6873 26736 6876
rect 26733 6872 26736 6873
rect 26762 6872 26765 6898
rect 29309 6872 29312 6898
rect 29338 6872 29341 6898
rect 24140 6844 24180 6858
rect 24319 6859 24348 6862
rect 24140 6838 24143 6844
rect 24319 6842 24325 6859
rect 24342 6858 24348 6859
rect 24571 6858 24574 6864
rect 24342 6844 24574 6858
rect 24342 6842 24348 6844
rect 24319 6839 24348 6842
rect 24571 6838 24574 6844
rect 24600 6838 24603 6864
rect 3036 6776 29992 6824
rect 14405 6736 14408 6762
rect 14434 6736 14437 6762
rect 22249 6757 22278 6760
rect 22249 6740 22255 6757
rect 22272 6756 22278 6757
rect 22639 6756 22642 6762
rect 22272 6742 22642 6756
rect 22272 6740 22278 6742
rect 22249 6737 22278 6740
rect 22639 6736 22642 6742
rect 22668 6736 22671 6762
rect 24847 6736 24850 6762
rect 24876 6756 24879 6762
rect 29033 6760 29036 6762
rect 25009 6757 25038 6760
rect 25009 6756 25015 6757
rect 24876 6742 25015 6756
rect 24876 6736 24879 6742
rect 25009 6740 25015 6742
rect 25032 6740 25038 6757
rect 25009 6737 25038 6740
rect 29011 6757 29036 6760
rect 29011 6740 29017 6757
rect 29034 6740 29036 6757
rect 29011 6737 29036 6740
rect 29033 6736 29036 6737
rect 29062 6736 29065 6762
rect 6079 6702 6082 6728
rect 6108 6722 6111 6728
rect 6108 6708 6976 6722
rect 6108 6702 6111 6708
rect 6217 6668 6220 6694
rect 6246 6668 6249 6694
rect 6962 6692 6976 6708
rect 6954 6689 6983 6692
rect 6954 6672 6960 6689
rect 6977 6672 6983 6689
rect 6954 6669 6983 6672
rect 10817 6668 10820 6694
rect 10846 6668 10849 6694
rect 10956 6689 10985 6692
rect 10956 6672 10962 6689
rect 10979 6688 10985 6689
rect 11139 6688 11142 6694
rect 10979 6674 11142 6688
rect 10979 6672 10985 6674
rect 10956 6669 10985 6672
rect 11139 6668 11142 6674
rect 11168 6668 11171 6694
rect 19282 6689 19311 6692
rect 19282 6672 19288 6689
rect 19305 6688 19311 6689
rect 20247 6688 20250 6694
rect 19305 6674 20250 6688
rect 19305 6672 19311 6674
rect 19282 6669 19311 6672
rect 20247 6668 20250 6674
rect 20276 6688 20279 6694
rect 20276 6674 21282 6688
rect 20276 6668 20279 6674
rect 6080 6655 6109 6658
rect 6080 6638 6086 6655
rect 6103 6654 6109 6655
rect 6226 6654 6240 6668
rect 21268 6660 21282 6674
rect 23237 6668 23240 6694
rect 23266 6688 23269 6694
rect 23973 6688 23976 6694
rect 23266 6674 23976 6688
rect 23266 6668 23269 6674
rect 23973 6668 23976 6674
rect 24002 6668 24005 6694
rect 27975 6668 27978 6694
rect 28004 6668 28007 6694
rect 6103 6640 6240 6654
rect 6816 6655 6845 6658
rect 6103 6638 6109 6640
rect 6080 6635 6109 6638
rect 6816 6638 6822 6655
rect 6839 6638 6845 6655
rect 6816 6635 6845 6638
rect 6862 6655 6891 6658
rect 6862 6638 6868 6655
rect 6885 6654 6891 6655
rect 7781 6654 7784 6660
rect 6885 6640 7784 6654
rect 6885 6638 6891 6640
rect 6862 6635 6891 6638
rect 5942 6621 5971 6624
rect 5942 6604 5948 6621
rect 5965 6620 5971 6621
rect 6217 6620 6220 6626
rect 5965 6606 6220 6620
rect 5965 6604 5971 6606
rect 5942 6601 5971 6604
rect 6217 6600 6220 6606
rect 6246 6600 6249 6626
rect 6824 6620 6838 6635
rect 7781 6634 7784 6640
rect 7810 6634 7813 6660
rect 13623 6634 13626 6660
rect 13652 6654 13655 6660
rect 13716 6655 13745 6658
rect 13716 6654 13722 6655
rect 13652 6640 13722 6654
rect 13652 6634 13655 6640
rect 13716 6638 13722 6640
rect 13739 6638 13745 6655
rect 13716 6635 13745 6638
rect 13761 6634 13764 6660
rect 13790 6654 13793 6660
rect 13844 6655 13873 6658
rect 13844 6654 13850 6655
rect 13790 6640 13850 6654
rect 13790 6634 13793 6640
rect 13844 6638 13850 6640
rect 13867 6638 13873 6655
rect 13844 6635 13873 6638
rect 17855 6634 17858 6660
rect 17884 6634 17887 6660
rect 17948 6655 17977 6658
rect 17948 6638 17954 6655
rect 17971 6654 17977 6655
rect 18085 6654 18088 6660
rect 17971 6640 18088 6654
rect 17971 6638 17977 6640
rect 17948 6635 17977 6638
rect 6907 6620 6910 6626
rect 6824 6606 6910 6620
rect 6907 6600 6910 6606
rect 6936 6600 6939 6626
rect 11001 6600 11004 6626
rect 11030 6620 11033 6626
rect 11030 6606 11201 6620
rect 11030 6600 11033 6606
rect 11829 6600 11832 6626
rect 11858 6600 11861 6626
rect 16107 6600 16110 6626
rect 16136 6620 16139 6626
rect 17956 6620 17970 6635
rect 18085 6634 18088 6640
rect 18114 6634 18117 6660
rect 18959 6634 18962 6660
rect 18988 6634 18991 6660
rect 19143 6634 19146 6660
rect 19172 6634 19175 6660
rect 19327 6634 19330 6660
rect 19356 6654 19359 6660
rect 19558 6655 19587 6658
rect 19558 6654 19564 6655
rect 19356 6640 19564 6654
rect 19356 6634 19359 6640
rect 19558 6638 19564 6640
rect 19581 6638 19587 6655
rect 19558 6635 19587 6638
rect 19788 6655 19817 6658
rect 19788 6638 19794 6655
rect 19811 6638 19817 6655
rect 19788 6635 19817 6638
rect 16136 6606 17970 6620
rect 19152 6620 19166 6634
rect 19796 6620 19810 6635
rect 21075 6634 21078 6660
rect 21104 6654 21107 6660
rect 21214 6655 21243 6658
rect 21214 6654 21220 6655
rect 21104 6640 21220 6654
rect 21104 6634 21107 6640
rect 21214 6638 21220 6640
rect 21237 6638 21243 6655
rect 21214 6635 21243 6638
rect 21259 6634 21262 6660
rect 21288 6634 21291 6660
rect 21351 6634 21354 6660
rect 21380 6658 21383 6660
rect 21380 6655 21398 6658
rect 21392 6638 21398 6655
rect 21380 6635 21398 6638
rect 21380 6634 21383 6635
rect 24111 6634 24114 6660
rect 24140 6658 24143 6660
rect 24140 6655 24158 6658
rect 24152 6638 24158 6655
rect 24140 6635 24158 6638
rect 28137 6655 28166 6658
rect 28137 6638 28143 6655
rect 28160 6654 28166 6655
rect 28389 6654 28392 6660
rect 28160 6640 28392 6654
rect 28160 6638 28166 6640
rect 28137 6635 28166 6638
rect 24140 6634 24143 6635
rect 28389 6634 28392 6640
rect 28418 6634 28421 6660
rect 19152 6606 19810 6620
rect 19926 6621 19955 6624
rect 16136 6600 16139 6606
rect 19926 6604 19932 6621
rect 19949 6620 19955 6621
rect 21121 6620 21124 6626
rect 19949 6606 21124 6620
rect 19949 6604 19955 6606
rect 19926 6601 19955 6604
rect 21121 6600 21124 6606
rect 21150 6600 21153 6626
rect 21443 6624 21446 6626
rect 21425 6621 21446 6624
rect 21425 6604 21431 6621
rect 21425 6601 21446 6604
rect 21443 6600 21446 6601
rect 21472 6600 21475 6626
rect 24203 6624 24206 6626
rect 24185 6621 24206 6624
rect 24185 6604 24191 6621
rect 24185 6601 24206 6604
rect 24203 6600 24206 6601
rect 24232 6600 24235 6626
rect 28205 6624 28208 6626
rect 28187 6621 28208 6624
rect 28187 6604 28193 6621
rect 28187 6601 28208 6604
rect 28205 6600 28208 6601
rect 28234 6600 28237 6626
rect 5987 6566 5990 6592
rect 6016 6590 6019 6592
rect 6016 6567 6020 6590
rect 6034 6587 6063 6590
rect 6034 6570 6040 6587
rect 6057 6586 6063 6587
rect 6125 6586 6128 6592
rect 6057 6572 6128 6586
rect 6057 6570 6063 6572
rect 6034 6567 6063 6570
rect 6016 6566 6019 6567
rect 6125 6566 6128 6572
rect 6154 6566 6157 6592
rect 6723 6566 6726 6592
rect 6752 6586 6755 6592
rect 6816 6587 6845 6590
rect 6816 6586 6822 6587
rect 6752 6572 6822 6586
rect 6752 6566 6755 6572
rect 6816 6570 6822 6572
rect 6839 6570 6845 6587
rect 6816 6567 6845 6570
rect 17902 6587 17931 6590
rect 17902 6570 17908 6587
rect 17925 6586 17931 6587
rect 18131 6586 18134 6592
rect 17925 6572 18134 6586
rect 17925 6570 17931 6572
rect 17902 6567 17931 6570
rect 18131 6566 18134 6572
rect 18160 6566 18163 6592
rect 3036 6504 29992 6552
rect 6125 6464 6128 6490
rect 6154 6464 6157 6490
rect 22111 6485 22140 6488
rect 6548 6470 6930 6484
rect 6080 6451 6109 6454
rect 6080 6434 6086 6451
rect 6103 6450 6109 6451
rect 6217 6450 6220 6456
rect 6103 6436 6220 6450
rect 6103 6434 6109 6436
rect 6080 6431 6109 6434
rect 6217 6430 6220 6436
rect 6246 6450 6249 6456
rect 6493 6450 6496 6456
rect 6246 6436 6496 6450
rect 6246 6430 6249 6436
rect 6493 6430 6496 6436
rect 6522 6430 6525 6456
rect 6034 6417 6063 6420
rect 6034 6400 6040 6417
rect 6057 6416 6063 6417
rect 6171 6416 6174 6422
rect 6057 6402 6174 6416
rect 6057 6400 6063 6402
rect 6034 6397 6063 6400
rect 6171 6396 6174 6402
rect 6200 6396 6203 6422
rect 6264 6417 6293 6420
rect 6264 6400 6270 6417
rect 6287 6400 6293 6417
rect 6264 6397 6293 6400
rect 6079 6362 6082 6388
rect 6108 6382 6111 6388
rect 6272 6382 6286 6397
rect 6108 6368 6286 6382
rect 6108 6362 6111 6368
rect 5941 6328 5944 6354
rect 5970 6348 5973 6354
rect 6548 6348 6562 6470
rect 6723 6430 6726 6456
rect 6752 6430 6755 6456
rect 6916 6450 6930 6470
rect 22111 6468 22117 6485
rect 22134 6484 22140 6485
rect 22731 6484 22734 6490
rect 22134 6470 22734 6484
rect 22134 6468 22140 6470
rect 22111 6465 22140 6468
rect 22731 6464 22734 6470
rect 22760 6464 22763 6490
rect 24341 6464 24344 6490
rect 24370 6484 24373 6490
rect 24710 6485 24739 6488
rect 24370 6470 24640 6484
rect 24370 6464 24373 6470
rect 7597 6450 7600 6456
rect 6916 6436 6969 6450
rect 7337 6436 7600 6450
rect 7597 6430 7600 6436
rect 7626 6430 7629 6456
rect 15923 6430 15926 6456
rect 15952 6450 15955 6456
rect 16015 6450 16018 6456
rect 15952 6436 16018 6450
rect 15952 6430 15955 6436
rect 16015 6430 16018 6436
rect 16044 6450 16047 6456
rect 16062 6451 16091 6454
rect 16062 6450 16068 6451
rect 16044 6436 16068 6450
rect 16044 6430 16047 6436
rect 16062 6434 16068 6436
rect 16085 6434 16091 6451
rect 17258 6451 17287 6454
rect 17258 6450 17264 6451
rect 16062 6431 16091 6434
rect 16622 6436 17264 6450
rect 15969 6396 15972 6422
rect 15998 6396 16001 6422
rect 16107 6396 16110 6422
rect 16136 6396 16139 6422
rect 16622 6420 16636 6436
rect 17258 6434 17264 6436
rect 17281 6450 17287 6451
rect 17855 6450 17858 6456
rect 17281 6436 17858 6450
rect 17281 6434 17287 6436
rect 17258 6431 17287 6434
rect 17855 6430 17858 6436
rect 17884 6430 17887 6456
rect 19143 6450 19146 6456
rect 18324 6436 19146 6450
rect 16522 6417 16551 6420
rect 16522 6400 16528 6417
rect 16545 6400 16551 6417
rect 16522 6397 16551 6400
rect 16614 6417 16643 6420
rect 16614 6400 16620 6417
rect 16637 6400 16643 6417
rect 16614 6397 16643 6400
rect 6585 6362 6588 6388
rect 6614 6362 6617 6388
rect 7597 6362 7600 6388
rect 7626 6362 7629 6388
rect 16291 6382 16294 6388
rect 16116 6368 16294 6382
rect 16116 6352 16130 6368
rect 16291 6362 16294 6368
rect 16320 6382 16323 6388
rect 16530 6382 16544 6397
rect 17119 6396 17122 6422
rect 17148 6396 17151 6422
rect 17166 6417 17195 6420
rect 17166 6400 17172 6417
rect 17189 6400 17195 6417
rect 17166 6397 17195 6400
rect 16320 6368 16544 6382
rect 16320 6362 16323 6368
rect 17027 6362 17030 6388
rect 17056 6382 17059 6388
rect 17174 6382 17188 6397
rect 18131 6396 18134 6422
rect 18160 6396 18163 6422
rect 18324 6420 18338 6436
rect 19143 6430 19146 6436
rect 19172 6430 19175 6456
rect 19327 6450 19330 6456
rect 19198 6436 19330 6450
rect 18316 6417 18345 6420
rect 18316 6400 18322 6417
rect 18339 6400 18345 6417
rect 18316 6397 18345 6400
rect 18407 6396 18410 6422
rect 18436 6396 18439 6422
rect 19098 6417 19127 6420
rect 19098 6400 19104 6417
rect 19121 6416 19127 6417
rect 19198 6416 19212 6436
rect 19327 6430 19330 6436
rect 19356 6430 19359 6456
rect 19373 6430 19376 6456
rect 19402 6430 19405 6456
rect 20118 6436 20454 6450
rect 20118 6422 20132 6436
rect 19121 6402 19212 6416
rect 19236 6417 19265 6420
rect 19121 6400 19127 6402
rect 19098 6397 19127 6400
rect 19236 6400 19242 6417
rect 19259 6416 19265 6417
rect 20109 6416 20112 6422
rect 19259 6402 20112 6416
rect 19259 6400 19265 6402
rect 19236 6397 19265 6400
rect 17056 6368 17188 6382
rect 17056 6362 17059 6368
rect 18683 6362 18686 6388
rect 18712 6382 18715 6388
rect 19244 6382 19258 6397
rect 20109 6396 20112 6402
rect 20138 6396 20141 6422
rect 20201 6396 20204 6422
rect 20230 6396 20233 6422
rect 20440 6420 20454 6436
rect 20569 6430 20572 6456
rect 20598 6430 20601 6456
rect 21305 6454 21308 6456
rect 21287 6451 21308 6454
rect 21287 6434 21293 6451
rect 21287 6431 21308 6434
rect 21305 6430 21308 6431
rect 21334 6430 21337 6456
rect 23375 6454 23378 6456
rect 23357 6451 23378 6454
rect 23357 6434 23363 6451
rect 23357 6431 23378 6434
rect 23375 6430 23378 6431
rect 23404 6430 23407 6456
rect 24534 6454 24548 6470
rect 24526 6451 24555 6454
rect 24526 6434 24532 6451
rect 24549 6434 24555 6451
rect 24526 6431 24555 6434
rect 24571 6430 24574 6456
rect 24600 6430 24603 6456
rect 24626 6450 24640 6470
rect 24710 6468 24716 6485
rect 24733 6484 24739 6485
rect 24755 6484 24758 6490
rect 24733 6470 24758 6484
rect 24733 6468 24739 6470
rect 24710 6465 24739 6468
rect 24755 6464 24758 6470
rect 24784 6464 24787 6490
rect 25445 6450 25448 6456
rect 24626 6436 25448 6450
rect 25445 6430 25448 6436
rect 25474 6430 25477 6456
rect 28417 6451 28446 6454
rect 28417 6434 28423 6451
rect 28440 6450 28446 6451
rect 28481 6450 28484 6456
rect 28440 6436 28484 6450
rect 28440 6434 28446 6436
rect 28417 6431 28446 6434
rect 28481 6430 28484 6436
rect 28510 6430 28513 6456
rect 20432 6417 20461 6420
rect 20432 6400 20438 6417
rect 20455 6400 20461 6417
rect 20432 6397 20461 6400
rect 21075 6396 21078 6422
rect 21104 6396 21107 6422
rect 21237 6417 21266 6420
rect 21237 6400 21243 6417
rect 21260 6416 21266 6417
rect 21351 6416 21354 6422
rect 21260 6402 21354 6416
rect 21260 6400 21266 6402
rect 21237 6397 21266 6400
rect 21351 6396 21354 6402
rect 21380 6396 21383 6422
rect 23146 6417 23175 6420
rect 23146 6400 23152 6417
rect 23169 6416 23175 6417
rect 23191 6416 23194 6422
rect 23169 6402 23194 6416
rect 23169 6400 23175 6402
rect 23146 6397 23175 6400
rect 23191 6396 23194 6402
rect 23220 6396 23223 6422
rect 23307 6417 23336 6420
rect 23307 6400 23313 6417
rect 23330 6416 23336 6417
rect 23559 6416 23562 6422
rect 23330 6402 23562 6416
rect 23330 6400 23336 6402
rect 23307 6397 23336 6400
rect 23559 6396 23562 6402
rect 23588 6396 23591 6422
rect 24181 6417 24210 6420
rect 24181 6400 24187 6417
rect 24204 6416 24210 6417
rect 24434 6417 24463 6420
rect 24434 6416 24440 6417
rect 24204 6402 24440 6416
rect 24204 6400 24210 6402
rect 24181 6397 24210 6400
rect 24434 6400 24440 6402
rect 24457 6400 24463 6417
rect 24434 6397 24463 6400
rect 24618 6417 24647 6420
rect 24618 6400 24624 6417
rect 24641 6400 24647 6417
rect 24618 6397 24647 6400
rect 18712 6368 19258 6382
rect 18712 6362 18715 6368
rect 5970 6334 6562 6348
rect 16108 6349 16137 6352
rect 5970 6328 5973 6334
rect 16108 6332 16114 6349
rect 16131 6332 16137 6349
rect 16108 6329 16137 6332
rect 5987 6294 5990 6320
rect 6016 6314 6019 6320
rect 6218 6315 6247 6318
rect 6218 6314 6224 6315
rect 6016 6300 6224 6314
rect 6016 6294 6019 6300
rect 6218 6298 6224 6300
rect 6241 6298 6247 6315
rect 6218 6295 6247 6298
rect 6263 6294 6266 6320
rect 6292 6294 6295 6320
rect 16521 6294 16524 6320
rect 16550 6294 16553 6320
rect 22961 6294 22964 6320
rect 22990 6314 22993 6320
rect 24626 6314 24640 6397
rect 27975 6396 27978 6422
rect 28004 6416 28007 6422
rect 28205 6416 28208 6422
rect 28004 6402 28208 6416
rect 28004 6396 28007 6402
rect 28205 6396 28208 6402
rect 28234 6396 28237 6422
rect 28343 6396 28346 6422
rect 28372 6420 28375 6422
rect 28372 6417 28390 6420
rect 28384 6400 28390 6417
rect 28372 6397 28390 6400
rect 28372 6396 28375 6397
rect 29171 6362 29174 6388
rect 29200 6382 29203 6388
rect 29241 6383 29270 6386
rect 29241 6382 29247 6383
rect 29200 6368 29247 6382
rect 29200 6362 29203 6368
rect 29241 6366 29247 6368
rect 29264 6366 29270 6383
rect 29241 6363 29270 6366
rect 22990 6300 24640 6314
rect 22990 6294 22993 6300
rect 3036 6232 29992 6280
rect 5527 6212 5530 6218
rect 5490 6198 5530 6212
rect 5490 6148 5504 6198
rect 5527 6192 5530 6198
rect 5556 6212 5559 6218
rect 6585 6212 6588 6218
rect 5556 6198 6588 6212
rect 5556 6192 5559 6198
rect 6585 6192 6588 6198
rect 6614 6192 6617 6218
rect 6907 6192 6910 6218
rect 6936 6212 6939 6218
rect 6954 6213 6983 6216
rect 6954 6212 6960 6213
rect 6936 6198 6960 6212
rect 6936 6192 6939 6198
rect 6954 6196 6960 6198
rect 6977 6196 6983 6213
rect 6954 6193 6983 6196
rect 6125 6158 6128 6184
rect 6154 6178 6157 6184
rect 6154 6164 6562 6178
rect 6154 6158 6157 6164
rect 5482 6145 5511 6148
rect 5482 6128 5488 6145
rect 5505 6128 5511 6145
rect 5482 6125 5511 6128
rect 5620 6145 5649 6148
rect 5620 6128 5626 6145
rect 5643 6144 5649 6145
rect 6263 6144 6266 6150
rect 5643 6130 6266 6144
rect 5643 6128 5649 6130
rect 5620 6125 5649 6128
rect 6263 6124 6266 6130
rect 6292 6124 6295 6150
rect 5941 6056 5944 6082
rect 5970 6056 5973 6082
rect 6493 6056 6496 6082
rect 6522 6056 6525 6082
rect 6548 6076 6562 6164
rect 6769 6158 6772 6184
rect 6798 6178 6801 6184
rect 7643 6178 7646 6184
rect 6798 6164 7646 6178
rect 6798 6158 6801 6164
rect 7643 6158 7646 6164
rect 7672 6158 7675 6184
rect 6778 6114 6792 6158
rect 6862 6145 6891 6148
rect 6862 6128 6868 6145
rect 6885 6144 6891 6145
rect 7414 6145 7443 6148
rect 7414 6144 7420 6145
rect 6885 6130 7420 6144
rect 6885 6128 6891 6130
rect 6862 6125 6891 6128
rect 7414 6128 7420 6130
rect 7437 6128 7443 6145
rect 7597 6144 7600 6150
rect 7414 6125 7443 6128
rect 7560 6130 7600 6144
rect 6770 6111 6799 6114
rect 6770 6094 6776 6111
rect 6793 6094 6799 6111
rect 6770 6091 6799 6094
rect 6870 6076 6884 6125
rect 7560 6114 7574 6130
rect 7597 6124 7600 6130
rect 7626 6144 7629 6150
rect 8011 6144 8014 6150
rect 7626 6130 8014 6144
rect 7626 6124 7629 6130
rect 8011 6124 8014 6130
rect 8040 6124 8043 6150
rect 20202 6145 20231 6148
rect 20202 6128 20208 6145
rect 20225 6144 20231 6145
rect 21305 6144 21308 6150
rect 20225 6130 21308 6144
rect 20225 6128 20231 6130
rect 20202 6125 20231 6128
rect 21305 6124 21308 6130
rect 21334 6124 21337 6150
rect 6954 6111 6983 6114
rect 6954 6094 6960 6111
rect 6977 6110 6983 6111
rect 7552 6111 7581 6114
rect 7552 6110 7558 6111
rect 6977 6096 7558 6110
rect 6977 6094 6983 6096
rect 6954 6091 6983 6094
rect 7552 6094 7558 6096
rect 7575 6094 7581 6111
rect 7552 6091 7581 6094
rect 7781 6090 7784 6116
rect 7810 6090 7813 6116
rect 11047 6090 11050 6116
rect 11076 6110 11079 6116
rect 11204 6111 11233 6114
rect 11204 6110 11210 6111
rect 11076 6096 11210 6110
rect 11076 6090 11079 6096
rect 11204 6094 11210 6096
rect 11227 6094 11233 6111
rect 11204 6091 11233 6094
rect 19879 6090 19882 6116
rect 19908 6090 19911 6116
rect 19971 6090 19974 6116
rect 20000 6110 20003 6116
rect 20018 6111 20047 6114
rect 20018 6110 20024 6111
rect 20000 6096 20024 6110
rect 20000 6090 20003 6096
rect 20018 6094 20024 6096
rect 20041 6094 20047 6111
rect 20018 6091 20047 6094
rect 20110 6111 20139 6114
rect 20110 6094 20116 6111
rect 20133 6110 20139 6111
rect 20155 6110 20158 6116
rect 20133 6096 20158 6110
rect 20133 6094 20139 6096
rect 20110 6091 20139 6094
rect 20155 6090 20158 6096
rect 20184 6090 20187 6116
rect 6548 6062 6884 6076
rect 7414 6077 7443 6080
rect 7414 6060 7420 6077
rect 7437 6076 7443 6077
rect 7598 6077 7627 6080
rect 7437 6062 7574 6076
rect 7437 6060 7443 6062
rect 7414 6057 7443 6060
rect 6502 6042 6516 6056
rect 6816 6043 6845 6046
rect 6816 6042 6822 6043
rect 6502 6028 6822 6042
rect 6816 6026 6822 6028
rect 6839 6042 6845 6043
rect 7505 6042 7508 6048
rect 6839 6028 7508 6042
rect 6839 6026 6845 6028
rect 6816 6023 6845 6026
rect 7505 6022 7508 6028
rect 7534 6022 7537 6048
rect 7560 6042 7574 6062
rect 7598 6060 7604 6077
rect 7621 6076 7627 6077
rect 7643 6076 7646 6082
rect 7621 6062 7646 6076
rect 7621 6060 7627 6062
rect 7598 6057 7627 6060
rect 7643 6056 7646 6062
rect 7672 6056 7675 6082
rect 9253 6042 9256 6048
rect 7560 6028 9256 6042
rect 9253 6022 9256 6028
rect 9282 6022 9285 6048
rect 11255 6043 11284 6046
rect 11255 6026 11261 6043
rect 11278 6042 11284 6043
rect 11553 6042 11556 6048
rect 11278 6028 11556 6042
rect 11278 6026 11284 6028
rect 11255 6023 11284 6026
rect 11553 6022 11556 6028
rect 11582 6022 11585 6048
rect 3036 5960 29992 6008
rect 7505 5920 7508 5946
rect 7534 5940 7537 5946
rect 11048 5941 11077 5944
rect 7534 5926 9506 5940
rect 7534 5920 7537 5926
rect 9492 5912 9506 5926
rect 11048 5924 11054 5941
rect 11071 5940 11077 5941
rect 11093 5940 11096 5946
rect 11071 5926 11096 5940
rect 11071 5924 11077 5926
rect 11048 5921 11077 5924
rect 11093 5920 11096 5926
rect 11122 5920 11125 5946
rect 18545 5920 18548 5946
rect 18574 5920 18577 5946
rect 29333 5941 29362 5944
rect 29333 5924 29339 5941
rect 29356 5940 29362 5941
rect 29677 5940 29680 5946
rect 29356 5926 29680 5940
rect 29356 5924 29362 5926
rect 29333 5921 29362 5924
rect 29677 5920 29680 5926
rect 29706 5920 29709 5946
rect 7827 5906 7830 5912
rect 7698 5892 7830 5906
rect 7698 5876 7712 5892
rect 7827 5886 7830 5892
rect 7856 5906 7859 5912
rect 8241 5906 8244 5912
rect 7856 5892 8244 5906
rect 7856 5886 7859 5892
rect 8241 5886 8244 5892
rect 8270 5886 8273 5912
rect 9253 5886 9256 5912
rect 9282 5906 9285 5912
rect 9282 5892 9368 5906
rect 9282 5886 9285 5892
rect 7690 5873 7719 5876
rect 7690 5856 7696 5873
rect 7713 5856 7719 5873
rect 7690 5853 7719 5856
rect 7735 5852 7738 5878
rect 7764 5872 7767 5878
rect 7782 5873 7811 5876
rect 7782 5872 7788 5873
rect 7764 5858 7788 5872
rect 7764 5852 7767 5858
rect 7782 5856 7788 5858
rect 7805 5872 7811 5873
rect 8150 5873 8179 5876
rect 8150 5872 8156 5873
rect 7805 5858 8156 5872
rect 7805 5856 7811 5858
rect 7782 5853 7811 5856
rect 8150 5856 8156 5858
rect 8173 5856 8179 5873
rect 8150 5853 8179 5856
rect 9299 5852 9302 5878
rect 9328 5852 9331 5878
rect 9354 5876 9368 5892
rect 9483 5886 9486 5912
rect 9512 5886 9515 5912
rect 10266 5907 10295 5910
rect 10266 5890 10272 5907
rect 10289 5906 10295 5907
rect 10449 5906 10452 5912
rect 10289 5892 10452 5906
rect 10289 5890 10295 5892
rect 10266 5887 10295 5890
rect 10449 5886 10452 5892
rect 10478 5886 10481 5912
rect 10956 5907 10985 5910
rect 10956 5890 10962 5907
rect 10979 5906 10985 5907
rect 11829 5906 11832 5912
rect 10979 5892 11832 5906
rect 10979 5890 10985 5892
rect 10956 5887 10985 5890
rect 9347 5873 9376 5876
rect 9347 5856 9353 5873
rect 9370 5856 9376 5873
rect 9347 5853 9376 5856
rect 9437 5852 9440 5878
rect 9466 5852 9469 5878
rect 9529 5852 9532 5878
rect 9558 5876 9561 5878
rect 9558 5872 9562 5876
rect 9852 5873 9881 5876
rect 9558 5858 9580 5872
rect 9558 5853 9562 5858
rect 9852 5856 9858 5873
rect 9875 5856 9881 5873
rect 9852 5853 9881 5856
rect 9990 5873 10019 5876
rect 9990 5856 9996 5873
rect 10013 5856 10019 5873
rect 9990 5853 10019 5856
rect 9558 5852 9561 5853
rect 8103 5818 8106 5844
rect 8132 5818 8135 5844
rect 9622 5805 9651 5808
rect 9622 5788 9628 5805
rect 9645 5804 9651 5805
rect 9860 5804 9874 5853
rect 9645 5790 9874 5804
rect 9998 5804 10012 5853
rect 10127 5852 10130 5878
rect 10156 5852 10159 5878
rect 10173 5852 10176 5878
rect 10202 5852 10205 5878
rect 11094 5873 11123 5876
rect 11094 5856 11100 5873
rect 11117 5856 11123 5873
rect 11094 5853 11123 5856
rect 11001 5818 11004 5844
rect 11030 5838 11033 5844
rect 11102 5838 11116 5853
rect 11553 5852 11556 5878
rect 11582 5852 11585 5878
rect 11700 5842 11714 5892
rect 11829 5886 11832 5892
rect 11858 5886 11861 5912
rect 18085 5886 18088 5912
rect 18114 5906 18117 5912
rect 18554 5906 18568 5920
rect 18960 5907 18989 5910
rect 18114 5892 18752 5906
rect 18114 5886 18117 5892
rect 17027 5852 17030 5878
rect 17056 5872 17059 5878
rect 17074 5873 17103 5876
rect 17074 5872 17080 5873
rect 17056 5858 17080 5872
rect 17056 5852 17059 5858
rect 17074 5856 17080 5858
rect 17097 5856 17103 5873
rect 17074 5853 17103 5856
rect 17119 5852 17122 5878
rect 17148 5872 17151 5878
rect 17211 5872 17214 5878
rect 17148 5858 17214 5872
rect 17148 5852 17151 5858
rect 17211 5852 17214 5858
rect 17240 5852 17243 5878
rect 17350 5873 17379 5876
rect 17350 5856 17356 5873
rect 17373 5872 17379 5873
rect 18269 5872 18272 5878
rect 17373 5858 18272 5872
rect 17373 5856 17379 5858
rect 17350 5853 17379 5856
rect 18269 5852 18272 5858
rect 18298 5872 18301 5878
rect 18362 5873 18391 5876
rect 18362 5872 18368 5873
rect 18298 5858 18368 5872
rect 18298 5852 18301 5858
rect 18362 5856 18368 5858
rect 18385 5856 18391 5873
rect 18362 5853 18391 5856
rect 18499 5852 18502 5878
rect 18528 5872 18531 5878
rect 18738 5876 18752 5892
rect 18960 5890 18966 5907
rect 18983 5906 18989 5907
rect 19097 5906 19100 5912
rect 18983 5892 19100 5906
rect 18983 5890 18989 5892
rect 18960 5887 18989 5890
rect 19097 5886 19100 5892
rect 19126 5906 19129 5912
rect 20202 5907 20231 5910
rect 19126 5892 20086 5906
rect 19126 5886 19129 5892
rect 18546 5873 18575 5876
rect 18546 5872 18552 5873
rect 18528 5858 18552 5872
rect 18528 5852 18531 5858
rect 18546 5856 18552 5858
rect 18569 5856 18575 5873
rect 18546 5853 18575 5856
rect 18730 5873 18759 5876
rect 18730 5856 18736 5873
rect 18753 5856 18759 5873
rect 18730 5853 18759 5856
rect 19327 5852 19330 5878
rect 19356 5872 19359 5878
rect 19833 5872 19836 5878
rect 19356 5858 19836 5872
rect 19356 5852 19359 5858
rect 19833 5852 19836 5858
rect 19862 5852 19865 5878
rect 20072 5876 20086 5892
rect 20202 5890 20208 5907
rect 20225 5906 20231 5907
rect 20707 5906 20710 5912
rect 20225 5892 20710 5906
rect 20225 5890 20231 5892
rect 20202 5887 20231 5890
rect 20707 5886 20710 5892
rect 20736 5886 20739 5912
rect 26227 5886 26230 5912
rect 26256 5906 26259 5912
rect 26619 5907 26648 5910
rect 26619 5906 26625 5907
rect 26256 5892 26625 5906
rect 26256 5886 26259 5892
rect 26619 5890 26625 5892
rect 26642 5890 26648 5907
rect 26619 5887 26648 5890
rect 28509 5907 28538 5910
rect 28509 5890 28515 5907
rect 28532 5906 28538 5907
rect 28573 5906 28576 5912
rect 28532 5892 28576 5906
rect 28532 5890 28538 5892
rect 28509 5887 28538 5890
rect 28573 5886 28576 5892
rect 28602 5886 28605 5912
rect 20064 5873 20093 5876
rect 20064 5856 20070 5873
rect 20087 5856 20093 5873
rect 20064 5853 20093 5856
rect 24203 5852 24206 5878
rect 24232 5872 24235 5878
rect 26567 5873 26596 5876
rect 26567 5872 26573 5873
rect 24232 5858 26573 5872
rect 24232 5852 24235 5858
rect 26567 5856 26573 5858
rect 26590 5872 26596 5873
rect 28343 5872 28346 5878
rect 26590 5858 28346 5872
rect 26590 5856 26596 5858
rect 26567 5853 26596 5856
rect 28343 5852 28346 5858
rect 28372 5872 28375 5878
rect 28453 5873 28482 5876
rect 28453 5872 28459 5873
rect 28372 5858 28459 5872
rect 28372 5852 28375 5858
rect 28453 5856 28459 5858
rect 28476 5856 28482 5873
rect 28453 5853 28482 5856
rect 11600 5839 11629 5842
rect 11600 5838 11606 5839
rect 11030 5824 11606 5838
rect 11030 5818 11033 5824
rect 11600 5822 11606 5824
rect 11623 5822 11629 5839
rect 11600 5819 11629 5822
rect 11692 5839 11721 5842
rect 11692 5822 11698 5839
rect 11715 5822 11721 5839
rect 11692 5819 11721 5822
rect 20109 5818 20112 5844
rect 20138 5818 20141 5844
rect 26412 5839 26441 5842
rect 26412 5822 26418 5839
rect 26435 5822 26441 5839
rect 26412 5819 26441 5822
rect 28298 5839 28327 5842
rect 28298 5822 28304 5839
rect 28321 5822 28327 5839
rect 28298 5819 28327 5822
rect 10956 5805 10985 5808
rect 10956 5804 10962 5805
rect 9998 5790 10962 5804
rect 9645 5788 9651 5790
rect 9622 5785 9651 5788
rect 10956 5788 10962 5790
rect 10979 5788 10985 5805
rect 10956 5785 10985 5788
rect 7690 5771 7719 5774
rect 7690 5754 7696 5771
rect 7713 5770 7719 5771
rect 7873 5770 7876 5776
rect 7713 5756 7876 5770
rect 7713 5754 7719 5756
rect 7690 5751 7719 5754
rect 7873 5750 7876 5756
rect 7902 5750 7905 5776
rect 8288 5771 8317 5774
rect 8288 5754 8294 5771
rect 8311 5770 8317 5771
rect 9023 5770 9026 5776
rect 8311 5756 9026 5770
rect 8311 5754 8317 5756
rect 8288 5751 8317 5754
rect 9023 5750 9026 5756
rect 9052 5750 9055 5776
rect 11645 5750 11648 5776
rect 11674 5750 11677 5776
rect 15923 5750 15926 5776
rect 15952 5770 15955 5776
rect 17212 5771 17241 5774
rect 17212 5770 17218 5771
rect 15952 5756 17218 5770
rect 15952 5750 15955 5756
rect 17212 5754 17218 5756
rect 17235 5754 17241 5771
rect 26420 5770 26434 5819
rect 28205 5804 28208 5810
rect 27248 5790 28208 5804
rect 27248 5770 27262 5790
rect 28205 5784 28208 5790
rect 28234 5804 28237 5810
rect 28306 5804 28320 5819
rect 28234 5790 28320 5804
rect 28234 5784 28237 5790
rect 26420 5756 27262 5770
rect 17212 5751 17241 5754
rect 27285 5750 27288 5776
rect 27314 5770 27317 5776
rect 27447 5771 27476 5774
rect 27447 5770 27453 5771
rect 27314 5756 27453 5770
rect 27314 5750 27317 5756
rect 27447 5754 27453 5756
rect 27470 5754 27476 5771
rect 27447 5751 27476 5754
rect 3036 5688 29992 5736
rect 10127 5648 10130 5674
rect 10156 5668 10159 5674
rect 10266 5669 10295 5672
rect 10266 5668 10272 5669
rect 10156 5654 10272 5668
rect 10156 5648 10159 5654
rect 10266 5652 10272 5654
rect 10289 5652 10295 5669
rect 17948 5669 17977 5672
rect 17948 5668 17954 5669
rect 10266 5649 10295 5652
rect 17220 5654 17954 5668
rect 7828 5635 7857 5638
rect 7828 5618 7834 5635
rect 7851 5634 7857 5635
rect 7851 5620 9092 5634
rect 7851 5618 7857 5620
rect 7828 5615 7857 5618
rect 7873 5580 7876 5606
rect 7902 5580 7905 5606
rect 7827 5546 7830 5572
rect 7856 5546 7859 5572
rect 7919 5546 7922 5572
rect 7948 5546 7951 5572
rect 8011 5546 8014 5572
rect 8040 5546 8043 5572
rect 8518 5567 8547 5570
rect 8518 5566 8524 5567
rect 8273 5552 8524 5566
rect 7735 5512 7738 5538
rect 7764 5532 7767 5538
rect 8273 5532 8287 5552
rect 8518 5550 8524 5552
rect 8541 5550 8547 5567
rect 8518 5547 8547 5550
rect 8609 5546 8612 5572
rect 8638 5546 8641 5572
rect 8932 5567 8961 5570
rect 8932 5550 8938 5567
rect 8955 5566 8961 5567
rect 8977 5566 8980 5572
rect 8955 5552 8980 5566
rect 8955 5550 8961 5552
rect 8932 5547 8961 5550
rect 8977 5546 8980 5552
rect 9006 5546 9009 5572
rect 9023 5546 9026 5572
rect 9052 5546 9055 5572
rect 9078 5570 9092 5620
rect 16567 5614 16570 5640
rect 16596 5634 16599 5640
rect 16596 5620 17004 5634
rect 16596 5614 16599 5620
rect 9483 5580 9486 5606
rect 9512 5600 9515 5606
rect 10174 5601 10203 5604
rect 10174 5600 10180 5601
rect 9512 5586 10180 5600
rect 9512 5580 9515 5586
rect 10174 5584 10180 5586
rect 10197 5584 10203 5601
rect 10174 5581 10203 5584
rect 10312 5601 10341 5604
rect 10312 5584 10318 5601
rect 10335 5600 10341 5601
rect 11645 5600 11648 5606
rect 10335 5586 11648 5600
rect 10335 5584 10341 5586
rect 10312 5581 10341 5584
rect 11645 5580 11648 5586
rect 11674 5580 11677 5606
rect 16061 5600 16064 5606
rect 15702 5586 16064 5600
rect 9070 5567 9099 5570
rect 9070 5550 9076 5567
rect 9093 5550 9099 5567
rect 9070 5547 9099 5550
rect 10219 5546 10222 5572
rect 10248 5546 10251 5572
rect 15702 5570 15716 5586
rect 16061 5580 16064 5586
rect 16090 5580 16093 5606
rect 16521 5600 16524 5606
rect 16392 5586 16524 5600
rect 15694 5567 15723 5570
rect 15694 5550 15700 5567
rect 15717 5550 15723 5567
rect 15694 5547 15723 5550
rect 15740 5567 15769 5570
rect 15740 5550 15746 5567
rect 15763 5566 15769 5567
rect 16392 5566 16406 5586
rect 16521 5580 16524 5586
rect 16550 5600 16553 5606
rect 16990 5604 17004 5620
rect 16890 5601 16919 5604
rect 16890 5600 16896 5601
rect 16550 5586 16896 5600
rect 16550 5580 16553 5586
rect 16890 5584 16896 5586
rect 16913 5584 16919 5601
rect 16890 5581 16919 5584
rect 16982 5601 17011 5604
rect 16982 5584 16988 5601
rect 17005 5600 17011 5601
rect 17027 5600 17030 5606
rect 17005 5586 17030 5600
rect 17005 5584 17011 5586
rect 16982 5581 17011 5584
rect 17027 5580 17030 5586
rect 17056 5580 17059 5606
rect 15763 5552 16406 5566
rect 16844 5567 16873 5570
rect 15763 5550 15769 5552
rect 15740 5547 15769 5550
rect 16844 5550 16850 5567
rect 16867 5566 16873 5567
rect 17220 5566 17234 5654
rect 17948 5652 17954 5654
rect 17971 5652 17977 5669
rect 17948 5649 17977 5652
rect 16867 5552 17234 5566
rect 17258 5567 17287 5570
rect 16867 5550 16873 5552
rect 16844 5547 16873 5550
rect 17258 5550 17264 5567
rect 17281 5550 17287 5567
rect 17956 5566 17970 5649
rect 18683 5648 18686 5674
rect 18712 5648 18715 5674
rect 19833 5648 19836 5674
rect 19862 5648 19865 5674
rect 22271 5634 22274 5640
rect 22234 5620 22274 5634
rect 19971 5600 19974 5606
rect 19796 5586 19974 5600
rect 18499 5566 18502 5572
rect 17956 5552 18502 5566
rect 17258 5547 17287 5550
rect 7764 5518 8287 5532
rect 8702 5533 8731 5536
rect 7764 5512 7767 5518
rect 8702 5516 8708 5533
rect 8725 5532 8731 5533
rect 9437 5532 9440 5538
rect 8725 5518 9440 5532
rect 8725 5516 8731 5518
rect 8702 5513 8731 5516
rect 9437 5512 9440 5518
rect 9466 5512 9469 5538
rect 15233 5512 15236 5538
rect 15262 5532 15265 5538
rect 15832 5533 15861 5536
rect 15832 5532 15838 5533
rect 15262 5518 15838 5532
rect 15262 5512 15265 5518
rect 15832 5516 15838 5518
rect 15855 5516 15861 5533
rect 15832 5513 15861 5516
rect 17119 5512 17122 5538
rect 17148 5532 17151 5538
rect 17266 5532 17280 5547
rect 18499 5546 18502 5552
rect 18528 5546 18531 5572
rect 18545 5546 18548 5572
rect 18574 5546 18577 5572
rect 18592 5567 18621 5570
rect 18592 5550 18598 5567
rect 18615 5550 18621 5567
rect 18592 5547 18621 5550
rect 17395 5536 17398 5538
rect 17148 5518 17280 5532
rect 17148 5512 17151 5518
rect 17392 5513 17398 5536
rect 17395 5512 17398 5513
rect 17424 5512 17427 5538
rect 18269 5512 18272 5538
rect 18298 5532 18301 5538
rect 18600 5532 18614 5547
rect 19603 5546 19606 5572
rect 19632 5566 19635 5572
rect 19796 5570 19810 5586
rect 19971 5580 19974 5586
rect 20000 5580 20003 5606
rect 19788 5567 19817 5570
rect 19788 5566 19794 5567
rect 19632 5552 19794 5566
rect 19632 5546 19635 5552
rect 19788 5550 19794 5552
rect 19811 5550 19817 5567
rect 19788 5547 19817 5550
rect 19879 5546 19882 5572
rect 19908 5566 19911 5572
rect 20064 5567 20093 5570
rect 20064 5566 20070 5567
rect 19908 5552 20070 5566
rect 19908 5546 19911 5552
rect 20064 5550 20070 5552
rect 20087 5550 20093 5567
rect 20064 5547 20093 5550
rect 22133 5546 22136 5572
rect 22162 5546 22165 5572
rect 22234 5570 22248 5620
rect 22271 5614 22274 5620
rect 22300 5634 22303 5640
rect 25399 5634 25402 5640
rect 22300 5620 25402 5634
rect 22300 5614 22303 5620
rect 25399 5614 25402 5620
rect 25428 5614 25431 5640
rect 26918 5601 26947 5604
rect 26918 5584 26924 5601
rect 26941 5600 26947 5601
rect 27009 5600 27012 5606
rect 26941 5586 27012 5600
rect 26941 5584 26947 5586
rect 26918 5581 26947 5584
rect 27009 5580 27012 5586
rect 27038 5580 27041 5606
rect 22211 5567 22248 5570
rect 22211 5550 22217 5567
rect 22234 5552 22248 5567
rect 22234 5550 22240 5552
rect 22211 5547 22240 5550
rect 22271 5546 22274 5572
rect 22300 5570 22303 5572
rect 22300 5567 22321 5570
rect 22315 5550 22321 5567
rect 22300 5547 22321 5550
rect 22347 5567 22376 5570
rect 22347 5550 22353 5567
rect 22370 5550 22376 5567
rect 22446 5567 22475 5570
rect 22347 5547 22376 5550
rect 22395 5557 22424 5560
rect 22300 5546 22303 5547
rect 18298 5518 18614 5532
rect 18298 5512 18301 5518
rect 21949 5512 21952 5538
rect 21978 5532 21981 5538
rect 22355 5532 22369 5547
rect 22395 5540 22401 5557
rect 22418 5555 22424 5557
rect 22418 5540 22432 5555
rect 22446 5550 22452 5567
rect 22469 5566 22475 5567
rect 22685 5566 22688 5572
rect 22469 5552 22688 5566
rect 22469 5550 22475 5552
rect 22446 5547 22475 5550
rect 22685 5546 22688 5552
rect 22714 5566 22717 5572
rect 22714 5552 23582 5566
rect 22714 5546 22717 5552
rect 22395 5537 22432 5540
rect 21978 5518 22369 5532
rect 21978 5512 21981 5518
rect 22418 5504 22432 5537
rect 23568 5532 23582 5552
rect 25353 5546 25356 5572
rect 25382 5566 25385 5572
rect 26734 5567 26763 5570
rect 26734 5566 26740 5567
rect 25382 5552 26740 5566
rect 25382 5546 25385 5552
rect 26734 5550 26740 5552
rect 26757 5550 26763 5567
rect 26734 5547 26763 5550
rect 26872 5567 26901 5570
rect 26872 5550 26878 5567
rect 26895 5550 26901 5567
rect 26872 5547 26901 5550
rect 25675 5532 25678 5538
rect 23568 5518 25678 5532
rect 25675 5512 25678 5518
rect 25704 5532 25707 5538
rect 26825 5532 26828 5538
rect 25704 5518 26828 5532
rect 25704 5512 25707 5518
rect 26825 5512 26828 5518
rect 26854 5512 26857 5538
rect 26880 5532 26894 5547
rect 27101 5546 27104 5572
rect 27130 5566 27133 5572
rect 27194 5567 27223 5570
rect 27194 5566 27200 5567
rect 27130 5552 27200 5566
rect 27130 5546 27133 5552
rect 27194 5550 27200 5552
rect 27217 5550 27223 5567
rect 27194 5547 27223 5550
rect 27285 5546 27288 5572
rect 27314 5546 27317 5572
rect 27240 5533 27269 5536
rect 27240 5532 27246 5533
rect 26880 5518 27246 5532
rect 27240 5516 27246 5518
rect 27263 5516 27269 5533
rect 27240 5513 27269 5516
rect 9070 5499 9099 5502
rect 9070 5482 9076 5499
rect 9093 5498 9099 5499
rect 10173 5498 10176 5504
rect 9093 5484 10176 5498
rect 9093 5482 9099 5484
rect 9070 5479 9099 5482
rect 10173 5478 10176 5484
rect 10202 5478 10205 5504
rect 15693 5478 15696 5504
rect 15722 5478 15725 5504
rect 16981 5478 16984 5504
rect 17010 5478 17013 5504
rect 22317 5478 22320 5504
rect 22346 5498 22349 5504
rect 22364 5499 22393 5502
rect 22364 5498 22370 5499
rect 22346 5484 22370 5498
rect 22346 5478 22349 5484
rect 22364 5482 22370 5484
rect 22387 5482 22393 5499
rect 22364 5479 22393 5482
rect 22409 5478 22412 5504
rect 22438 5478 22441 5504
rect 3036 5416 29992 5464
rect 7828 5397 7857 5400
rect 7828 5380 7834 5397
rect 7851 5396 7857 5397
rect 8011 5396 8014 5402
rect 7851 5382 8014 5396
rect 7851 5380 7857 5382
rect 7828 5377 7857 5380
rect 8011 5376 8014 5382
rect 8040 5376 8043 5402
rect 9116 5397 9145 5400
rect 9116 5380 9122 5397
rect 9139 5396 9145 5397
rect 9529 5396 9532 5402
rect 9139 5382 9532 5396
rect 9139 5380 9145 5382
rect 9116 5377 9145 5380
rect 9529 5376 9532 5382
rect 9558 5376 9561 5402
rect 10128 5397 10157 5400
rect 10128 5380 10134 5397
rect 10151 5396 10157 5397
rect 11001 5396 11004 5402
rect 10151 5382 11004 5396
rect 10151 5380 10157 5382
rect 10128 5377 10157 5380
rect 11001 5376 11004 5382
rect 11030 5376 11033 5402
rect 15969 5376 15972 5402
rect 15998 5376 16001 5402
rect 16061 5376 16064 5402
rect 16090 5376 16093 5402
rect 17395 5376 17398 5402
rect 17424 5376 17427 5402
rect 22111 5397 22140 5400
rect 22111 5380 22117 5397
rect 22134 5396 22140 5397
rect 22271 5396 22274 5402
rect 22134 5382 22274 5396
rect 22134 5380 22140 5382
rect 22111 5377 22140 5380
rect 22271 5376 22274 5382
rect 22300 5376 22303 5402
rect 25353 5376 25356 5402
rect 25382 5376 25385 5402
rect 25445 5376 25448 5402
rect 25474 5396 25477 5402
rect 25474 5382 25575 5396
rect 25474 5376 25477 5382
rect 7735 5342 7738 5368
rect 7764 5362 7767 5368
rect 9538 5362 9552 5376
rect 15138 5363 15167 5366
rect 7764 5348 8954 5362
rect 9538 5348 10150 5362
rect 7764 5342 7767 5348
rect 7782 5329 7811 5332
rect 7782 5312 7788 5329
rect 7805 5328 7811 5329
rect 7919 5328 7922 5334
rect 7805 5314 7922 5328
rect 7805 5312 7811 5314
rect 7782 5309 7811 5312
rect 7919 5308 7922 5314
rect 7948 5308 7951 5334
rect 7974 5332 7988 5348
rect 7966 5329 7995 5332
rect 7966 5312 7972 5329
rect 7989 5312 7995 5329
rect 7966 5309 7995 5312
rect 8196 5329 8225 5332
rect 8196 5312 8202 5329
rect 8219 5312 8225 5329
rect 8196 5309 8225 5312
rect 7874 5295 7903 5298
rect 7874 5278 7880 5295
rect 7897 5278 7903 5295
rect 8204 5294 8218 5309
rect 8287 5308 8290 5334
rect 8316 5308 8319 5334
rect 8940 5332 8954 5348
rect 8932 5329 8961 5332
rect 8932 5312 8938 5329
rect 8955 5312 8961 5329
rect 8932 5309 8961 5312
rect 8979 5329 9008 5332
rect 8979 5312 8985 5329
rect 9002 5312 9008 5329
rect 8979 5309 9008 5312
rect 7874 5275 7903 5278
rect 7974 5280 8218 5294
rect 7882 5226 7896 5275
rect 7974 5264 7988 5280
rect 8241 5274 8244 5300
rect 8270 5294 8273 5300
rect 8986 5294 9000 5309
rect 9437 5308 9440 5334
rect 9466 5328 9469 5334
rect 10136 5332 10150 5348
rect 15138 5346 15144 5363
rect 15161 5362 15167 5363
rect 15693 5362 15696 5368
rect 15161 5348 15696 5362
rect 15161 5346 15167 5348
rect 15138 5343 15167 5346
rect 15693 5342 15696 5348
rect 15722 5342 15725 5368
rect 17119 5362 17122 5368
rect 15863 5348 17122 5362
rect 10036 5329 10065 5332
rect 10036 5328 10042 5329
rect 9466 5314 10042 5328
rect 9466 5308 9469 5314
rect 10036 5312 10042 5314
rect 10059 5312 10065 5329
rect 10036 5309 10065 5312
rect 10128 5329 10157 5332
rect 10128 5312 10134 5329
rect 10151 5312 10157 5329
rect 10128 5309 10157 5312
rect 13623 5308 13626 5334
rect 13652 5328 13655 5334
rect 15004 5329 15033 5332
rect 15004 5328 15010 5329
rect 13652 5314 15010 5328
rect 13652 5308 13655 5314
rect 15004 5312 15010 5314
rect 15027 5328 15033 5329
rect 15863 5328 15877 5348
rect 17119 5342 17122 5348
rect 17148 5342 17151 5368
rect 20109 5362 20112 5368
rect 17450 5348 20112 5362
rect 15027 5314 15877 5328
rect 15027 5312 15033 5314
rect 15004 5309 15033 5312
rect 15923 5308 15926 5334
rect 15952 5308 15955 5334
rect 16107 5308 16110 5334
rect 16136 5308 16139 5334
rect 16981 5308 16984 5334
rect 17010 5328 17013 5334
rect 17450 5332 17464 5348
rect 20109 5342 20112 5348
rect 20138 5342 20141 5368
rect 20294 5363 20323 5366
rect 20294 5346 20300 5363
rect 20317 5362 20323 5363
rect 20845 5362 20848 5368
rect 20317 5348 20848 5362
rect 20317 5346 20323 5348
rect 20294 5343 20323 5346
rect 20845 5342 20848 5348
rect 20874 5342 20877 5368
rect 21305 5366 21308 5368
rect 21287 5363 21308 5366
rect 21287 5346 21293 5363
rect 21287 5343 21308 5346
rect 21305 5342 21308 5343
rect 21334 5342 21337 5368
rect 23375 5342 23378 5368
rect 23404 5362 23407 5368
rect 23997 5363 24026 5366
rect 23997 5362 24003 5363
rect 23404 5348 24003 5362
rect 23404 5342 23407 5348
rect 23997 5346 24003 5348
rect 24020 5346 24026 5363
rect 23997 5343 24026 5346
rect 25561 5343 25575 5382
rect 25560 5340 25589 5343
rect 17350 5329 17379 5332
rect 17350 5328 17356 5329
rect 17010 5314 17356 5328
rect 17010 5308 17013 5314
rect 17350 5312 17356 5314
rect 17373 5312 17379 5329
rect 17350 5309 17379 5312
rect 17442 5329 17471 5332
rect 17442 5312 17448 5329
rect 17465 5312 17471 5329
rect 17442 5309 17471 5312
rect 18269 5308 18272 5334
rect 18298 5328 18301 5334
rect 18362 5329 18391 5332
rect 18362 5328 18368 5329
rect 18298 5314 18368 5328
rect 18298 5308 18301 5314
rect 18362 5312 18368 5314
rect 18385 5312 18391 5329
rect 18362 5309 18391 5312
rect 18959 5308 18962 5334
rect 18988 5328 18991 5334
rect 19926 5329 19955 5332
rect 19926 5328 19932 5329
rect 18988 5314 19932 5328
rect 18988 5308 18991 5314
rect 19926 5312 19932 5314
rect 19949 5312 19955 5329
rect 19926 5309 19955 5312
rect 20155 5308 20158 5334
rect 20184 5308 20187 5334
rect 21075 5308 21078 5334
rect 21104 5308 21107 5334
rect 21237 5329 21266 5332
rect 21237 5312 21243 5329
rect 21260 5328 21266 5329
rect 21351 5328 21354 5334
rect 21260 5314 21354 5328
rect 21260 5312 21266 5314
rect 21237 5309 21266 5312
rect 21351 5308 21354 5314
rect 21380 5308 21383 5334
rect 23790 5329 23819 5332
rect 23790 5312 23796 5329
rect 23813 5328 23819 5329
rect 23835 5328 23838 5334
rect 23813 5314 23838 5328
rect 23813 5312 23819 5314
rect 23790 5309 23819 5312
rect 23835 5308 23838 5314
rect 23864 5308 23867 5334
rect 23951 5329 23980 5332
rect 23951 5312 23957 5329
rect 23974 5328 23980 5329
rect 24203 5328 24206 5334
rect 23974 5314 24206 5328
rect 23974 5312 23980 5314
rect 23951 5309 23980 5312
rect 24203 5308 24206 5314
rect 24232 5308 24235 5334
rect 25353 5308 25356 5334
rect 25382 5308 25385 5334
rect 25399 5308 25402 5334
rect 25428 5332 25431 5334
rect 25428 5329 25440 5332
rect 25434 5312 25440 5329
rect 25505 5329 25534 5332
rect 25505 5328 25511 5329
rect 25428 5309 25440 5312
rect 25500 5312 25511 5328
rect 25528 5312 25534 5329
rect 25560 5323 25566 5340
rect 25583 5323 25589 5340
rect 25675 5332 25678 5334
rect 25560 5320 25589 5323
rect 25615 5329 25644 5332
rect 25500 5309 25534 5312
rect 25615 5312 25621 5329
rect 25638 5328 25644 5329
rect 25666 5329 25678 5332
rect 25638 5312 25652 5328
rect 25615 5309 25652 5312
rect 25666 5312 25672 5329
rect 25666 5309 25678 5312
rect 25428 5308 25431 5309
rect 8270 5280 9000 5294
rect 8270 5274 8273 5280
rect 16015 5274 16018 5300
rect 16044 5274 16047 5300
rect 7966 5261 7995 5264
rect 7966 5244 7972 5261
rect 7989 5244 7995 5261
rect 7966 5241 7995 5244
rect 8196 5261 8225 5264
rect 8196 5244 8202 5261
rect 8219 5260 8225 5261
rect 10219 5260 10222 5266
rect 8219 5246 10222 5260
rect 8219 5244 8225 5246
rect 8196 5241 8225 5244
rect 10219 5240 10222 5246
rect 10248 5240 10251 5266
rect 15694 5261 15723 5264
rect 15694 5244 15700 5261
rect 15717 5260 15723 5261
rect 16116 5260 16130 5308
rect 18315 5294 18318 5300
rect 15717 5246 16130 5260
rect 16990 5280 18318 5294
rect 15717 5244 15723 5246
rect 15694 5241 15723 5244
rect 8287 5226 8290 5232
rect 7882 5212 8290 5226
rect 8287 5206 8290 5212
rect 8316 5226 8319 5232
rect 8609 5226 8612 5232
rect 8316 5212 8612 5226
rect 8316 5206 8319 5212
rect 8609 5206 8612 5212
rect 8638 5206 8641 5232
rect 16015 5206 16018 5232
rect 16044 5226 16047 5232
rect 16990 5226 17004 5280
rect 18315 5274 18318 5280
rect 18344 5274 18347 5300
rect 18454 5295 18483 5298
rect 18454 5278 18460 5295
rect 18477 5278 18483 5295
rect 18454 5275 18483 5278
rect 24825 5295 24854 5298
rect 24825 5278 24831 5295
rect 24848 5294 24854 5295
rect 25500 5294 25514 5309
rect 24848 5280 25514 5294
rect 24848 5278 24854 5280
rect 24825 5275 24854 5278
rect 17027 5240 17030 5266
rect 17056 5260 17059 5266
rect 18462 5260 18476 5275
rect 25638 5266 25652 5309
rect 25675 5308 25678 5309
rect 25704 5308 25707 5334
rect 17056 5246 18476 5260
rect 17056 5240 17059 5246
rect 25629 5240 25632 5266
rect 25658 5240 25661 5266
rect 16044 5212 17004 5226
rect 18408 5227 18437 5230
rect 16044 5206 16047 5212
rect 18408 5210 18414 5227
rect 18431 5226 18437 5227
rect 18637 5226 18640 5232
rect 18431 5212 18640 5226
rect 18431 5210 18437 5212
rect 18408 5207 18437 5210
rect 18637 5206 18640 5212
rect 18666 5206 18669 5232
rect 20845 5206 20848 5232
rect 20874 5226 20877 5232
rect 23375 5226 23378 5232
rect 20874 5212 23378 5226
rect 20874 5206 20877 5212
rect 23375 5206 23378 5212
rect 23404 5206 23407 5232
rect 3036 5144 29992 5192
rect 8173 5125 8202 5128
rect 8173 5108 8179 5125
rect 8196 5124 8202 5125
rect 8287 5124 8290 5130
rect 8196 5110 8290 5124
rect 8196 5108 8202 5110
rect 8173 5105 8202 5108
rect 8287 5104 8290 5110
rect 8316 5104 8319 5130
rect 22133 5104 22136 5130
rect 22162 5124 22165 5130
rect 22249 5125 22278 5128
rect 22249 5124 22255 5125
rect 22162 5110 22255 5124
rect 22162 5104 22165 5110
rect 22249 5108 22255 5110
rect 22272 5108 22278 5125
rect 22249 5105 22278 5108
rect 25009 5125 25038 5128
rect 25009 5108 25015 5125
rect 25032 5124 25038 5125
rect 25353 5124 25356 5130
rect 25032 5110 25356 5124
rect 25032 5108 25038 5110
rect 25009 5105 25038 5108
rect 25353 5104 25356 5110
rect 25382 5104 25385 5130
rect 18269 5036 18272 5062
rect 18298 5056 18301 5062
rect 18546 5057 18575 5060
rect 18546 5056 18552 5057
rect 18298 5042 18552 5056
rect 18298 5036 18301 5042
rect 18546 5040 18552 5042
rect 18569 5040 18575 5057
rect 18959 5056 18962 5062
rect 18546 5037 18575 5040
rect 18600 5042 18962 5056
rect 7827 5002 7830 5028
rect 7856 5022 7859 5028
rect 8122 5023 8151 5026
rect 8122 5022 8128 5023
rect 7856 5008 8128 5022
rect 7856 5002 7859 5008
rect 8122 5006 8128 5008
rect 8145 5022 8151 5023
rect 8241 5022 8244 5028
rect 8145 5008 8244 5022
rect 8145 5006 8151 5008
rect 8122 5003 8151 5006
rect 8241 5002 8244 5008
rect 8270 5002 8273 5028
rect 18454 5023 18483 5026
rect 18454 5006 18460 5023
rect 18477 5022 18483 5023
rect 18600 5022 18614 5042
rect 18959 5036 18962 5042
rect 18988 5056 18991 5062
rect 19742 5057 19771 5060
rect 19742 5056 19748 5057
rect 18988 5042 19748 5056
rect 18988 5036 18991 5042
rect 19742 5040 19748 5042
rect 19765 5040 19771 5057
rect 19742 5037 19771 5040
rect 21075 5036 21078 5062
rect 21104 5056 21107 5062
rect 21214 5057 21243 5060
rect 21214 5056 21220 5057
rect 21104 5042 21220 5056
rect 21104 5036 21107 5042
rect 21214 5040 21220 5042
rect 21237 5040 21243 5057
rect 21214 5037 21243 5040
rect 23835 5036 23838 5062
rect 23864 5056 23867 5062
rect 23974 5057 24003 5060
rect 23974 5056 23980 5057
rect 23864 5042 23980 5056
rect 23864 5036 23867 5042
rect 23974 5040 23980 5042
rect 23997 5040 24003 5057
rect 23974 5037 24003 5040
rect 18477 5008 18614 5022
rect 18477 5006 18483 5008
rect 18454 5003 18483 5006
rect 18637 5002 18640 5028
rect 18666 5002 18669 5028
rect 19603 5002 19606 5028
rect 19632 5002 19635 5028
rect 19879 5002 19882 5028
rect 19908 5022 19911 5028
rect 19926 5023 19955 5026
rect 19926 5022 19932 5023
rect 19908 5008 19932 5022
rect 19908 5002 19911 5008
rect 19926 5006 19932 5008
rect 19949 5006 19955 5023
rect 19926 5003 19955 5006
rect 21351 5002 21354 5028
rect 21380 5026 21383 5028
rect 21380 5023 21398 5026
rect 21392 5006 21398 5023
rect 21380 5003 21398 5006
rect 24135 5023 24164 5026
rect 24135 5006 24141 5023
rect 24158 5022 24164 5023
rect 24249 5022 24252 5028
rect 24158 5008 24252 5022
rect 24158 5006 24164 5008
rect 24135 5003 24164 5006
rect 21380 5002 21383 5003
rect 24249 5002 24252 5008
rect 24278 5002 24281 5028
rect 21443 4992 21446 4994
rect 21425 4989 21446 4992
rect 21425 4972 21431 4989
rect 21425 4969 21446 4972
rect 21443 4968 21446 4969
rect 21472 4968 21475 4994
rect 24203 4992 24206 4994
rect 24185 4989 24206 4992
rect 24185 4972 24191 4989
rect 24185 4969 24206 4972
rect 24203 4968 24206 4969
rect 24232 4968 24235 4994
rect 18453 4934 18456 4960
rect 18482 4954 18485 4960
rect 18500 4955 18529 4958
rect 18500 4954 18506 4955
rect 18482 4940 18506 4954
rect 18482 4934 18485 4940
rect 18500 4938 18506 4940
rect 18523 4938 18529 4955
rect 18500 4935 18529 4938
rect 18591 4934 18594 4960
rect 18620 4934 18623 4960
rect 3036 4872 29992 4920
rect 15969 4832 15972 4858
rect 15998 4852 16001 4858
rect 16522 4853 16551 4856
rect 16522 4852 16528 4853
rect 15998 4838 16528 4852
rect 15998 4832 16001 4838
rect 16522 4836 16528 4838
rect 16545 4836 16551 4853
rect 16522 4833 16551 4836
rect 15923 4798 15926 4824
rect 15952 4818 15955 4824
rect 16430 4819 16459 4822
rect 16430 4818 16436 4819
rect 15952 4804 16436 4818
rect 15952 4798 15955 4804
rect 16430 4802 16436 4804
rect 16453 4802 16459 4819
rect 16530 4818 16544 4833
rect 18315 4832 18318 4858
rect 18344 4852 18347 4858
rect 19098 4853 19127 4856
rect 19098 4852 19104 4853
rect 18344 4838 19104 4852
rect 18344 4832 18347 4838
rect 19098 4836 19104 4838
rect 19121 4836 19127 4853
rect 19098 4833 19127 4836
rect 17166 4819 17195 4822
rect 17166 4818 17172 4819
rect 16530 4804 17172 4818
rect 16430 4799 16459 4802
rect 17166 4802 17172 4804
rect 17189 4818 17195 4819
rect 17257 4818 17260 4824
rect 17189 4804 17260 4818
rect 17189 4802 17195 4804
rect 17166 4799 17195 4802
rect 17257 4798 17260 4804
rect 17286 4798 17289 4824
rect 18542 4819 18571 4822
rect 18542 4802 18548 4819
rect 18565 4818 18571 4819
rect 18591 4818 18594 4824
rect 18565 4804 18594 4818
rect 18565 4802 18571 4804
rect 18542 4799 18571 4802
rect 18591 4798 18594 4804
rect 18620 4798 18623 4824
rect 16568 4785 16597 4788
rect 16568 4768 16574 4785
rect 16591 4784 16597 4785
rect 17027 4784 17030 4790
rect 16591 4770 17030 4784
rect 16591 4768 16597 4770
rect 16568 4765 16597 4768
rect 17027 4764 17030 4770
rect 17056 4764 17059 4790
rect 17074 4785 17103 4788
rect 17074 4768 17080 4785
rect 17097 4768 17103 4785
rect 17074 4765 17103 4768
rect 16430 4717 16459 4720
rect 16430 4700 16436 4717
rect 16453 4716 16459 4717
rect 17082 4716 17096 4765
rect 17211 4764 17214 4790
rect 17240 4764 17243 4790
rect 18453 4764 18456 4790
rect 18482 4784 18485 4790
rect 19106 4784 19120 4833
rect 19603 4798 19606 4824
rect 19632 4818 19635 4824
rect 19632 4804 20178 4818
rect 19632 4798 19635 4804
rect 19834 4785 19863 4788
rect 19834 4784 19840 4785
rect 18482 4770 18982 4784
rect 19106 4770 19840 4784
rect 18482 4764 18485 4770
rect 17119 4730 17122 4756
rect 17148 4750 17151 4756
rect 18408 4751 18437 4754
rect 18408 4750 18414 4751
rect 17148 4736 18414 4750
rect 17148 4730 17151 4736
rect 18408 4734 18414 4736
rect 18431 4734 18437 4751
rect 18968 4750 18982 4770
rect 19834 4768 19840 4770
rect 19857 4784 19863 4785
rect 19879 4784 19882 4790
rect 19857 4770 19882 4784
rect 19857 4768 19863 4770
rect 19834 4765 19863 4768
rect 19879 4764 19882 4770
rect 19908 4764 19911 4790
rect 20164 4788 20178 4804
rect 21121 4798 21124 4824
rect 21150 4818 21153 4824
rect 21283 4819 21312 4822
rect 21283 4818 21289 4819
rect 21150 4804 21289 4818
rect 21150 4798 21153 4804
rect 21283 4802 21289 4804
rect 21306 4802 21312 4819
rect 21283 4799 21312 4802
rect 22111 4819 22140 4822
rect 22111 4802 22117 4819
rect 22134 4818 22140 4819
rect 22409 4818 22412 4824
rect 22134 4804 22412 4818
rect 22134 4802 22140 4804
rect 22111 4799 22140 4802
rect 22409 4798 22412 4804
rect 22438 4798 22441 4824
rect 20156 4785 20185 4788
rect 20156 4768 20162 4785
rect 20179 4768 20185 4785
rect 20156 4765 20185 4768
rect 21075 4764 21078 4790
rect 21104 4764 21107 4790
rect 21237 4785 21266 4788
rect 21237 4768 21243 4785
rect 21260 4784 21266 4785
rect 21351 4784 21354 4790
rect 21260 4770 21354 4784
rect 21260 4768 21266 4770
rect 21237 4765 21266 4768
rect 21351 4764 21354 4770
rect 21380 4764 21383 4790
rect 19972 4751 20001 4754
rect 19972 4750 19978 4751
rect 18968 4736 19978 4750
rect 18408 4731 18437 4734
rect 19972 4734 19978 4736
rect 19995 4734 20001 4751
rect 19972 4731 20001 4734
rect 16453 4702 17096 4716
rect 16453 4700 16459 4702
rect 16430 4697 16459 4700
rect 17073 4662 17076 4688
rect 17102 4662 17105 4688
rect 3036 4600 29992 4648
rect 17119 4580 17122 4586
rect 16576 4566 17122 4580
rect 16576 4516 16590 4566
rect 17119 4560 17122 4566
rect 17148 4560 17151 4586
rect 17257 4560 17260 4586
rect 17286 4580 17289 4586
rect 19603 4580 19606 4586
rect 17286 4566 19606 4580
rect 17286 4560 17289 4566
rect 19603 4560 19606 4566
rect 19632 4560 19635 4586
rect 25101 4581 25130 4584
rect 25101 4564 25107 4581
rect 25124 4580 25130 4581
rect 25629 4580 25632 4586
rect 25124 4566 25632 4580
rect 25124 4564 25130 4566
rect 25101 4561 25130 4564
rect 25629 4560 25632 4566
rect 25658 4560 25661 4586
rect 16568 4513 16597 4516
rect 16568 4496 16574 4513
rect 16591 4496 16597 4513
rect 16568 4493 16597 4496
rect 23835 4492 23838 4518
rect 23864 4512 23867 4518
rect 24066 4513 24095 4516
rect 24066 4512 24072 4513
rect 23864 4498 24072 4512
rect 23864 4492 23867 4498
rect 24066 4496 24072 4498
rect 24089 4496 24095 4513
rect 24066 4493 24095 4496
rect 16702 4479 16731 4482
rect 16702 4462 16708 4479
rect 16725 4478 16731 4479
rect 17073 4478 17076 4484
rect 16725 4464 17076 4478
rect 16725 4462 16731 4464
rect 16702 4459 16731 4462
rect 17073 4458 17076 4464
rect 17102 4458 17105 4484
rect 24203 4458 24206 4484
rect 24232 4482 24235 4484
rect 24232 4479 24250 4482
rect 24244 4462 24250 4479
rect 25951 4478 25954 4484
rect 24232 4459 24250 4462
rect 24350 4464 25954 4478
rect 24232 4458 24235 4459
rect 21121 4424 21124 4450
rect 21150 4444 21153 4450
rect 24273 4445 24302 4448
rect 24273 4444 24279 4445
rect 21150 4430 24279 4444
rect 21150 4424 21153 4430
rect 24273 4428 24279 4430
rect 24296 4444 24302 4445
rect 24350 4444 24364 4464
rect 25951 4458 25954 4464
rect 25980 4458 25983 4484
rect 24296 4430 24364 4444
rect 24296 4428 24302 4430
rect 24273 4425 24302 4428
rect 3036 4328 29992 4376
rect 3036 4056 29992 4104
rect 18637 3948 18640 3974
rect 18666 3948 18669 3974
rect 19098 3969 19127 3972
rect 19098 3952 19104 3969
rect 19121 3968 19127 3969
rect 19189 3968 19192 3974
rect 19121 3954 19192 3968
rect 19121 3952 19127 3954
rect 19098 3949 19127 3952
rect 19189 3948 19192 3954
rect 19218 3948 19221 3974
rect 18775 3914 18778 3940
rect 18804 3934 18807 3940
rect 20385 3934 20388 3940
rect 18804 3920 20388 3934
rect 18804 3914 18807 3920
rect 20385 3914 20388 3920
rect 20414 3914 20417 3940
rect 3036 3784 29992 3832
rect 3036 3512 29992 3560
rect 3036 3240 29992 3288
rect 16291 650 16294 676
rect 16320 670 16323 676
rect 16705 670 16708 676
rect 16320 656 16708 670
rect 16320 650 16323 656
rect 16705 650 16708 656
rect 16734 650 16737 676
<< via1 >>
rect 15880 29788 15906 29814
rect 16248 29686 16274 29712
rect 10268 29571 10294 29576
rect 10268 29554 10272 29571
rect 10272 29554 10289 29571
rect 10289 29554 10294 29571
rect 10268 29550 10294 29554
rect 15420 29550 15446 29576
rect 10360 29482 10386 29508
rect 10498 29482 10524 29508
rect 11372 29482 11398 29508
rect 12292 29482 12318 29508
rect 16340 29516 16366 29542
rect 8704 29448 8730 29474
rect 10544 29414 10570 29440
rect 11878 29448 11904 29474
rect 12338 29448 12364 29474
rect 15696 29469 15722 29474
rect 15696 29452 15700 29469
rect 15700 29452 15717 29469
rect 15717 29452 15722 29469
rect 15696 29448 15722 29452
rect 16202 29482 16228 29508
rect 12108 29435 12134 29440
rect 12108 29418 12112 29435
rect 12112 29418 12129 29435
rect 12129 29418 12134 29435
rect 12108 29414 12134 29418
rect 15788 29435 15814 29440
rect 15788 29418 15792 29435
rect 15792 29418 15809 29435
rect 15809 29418 15814 29435
rect 15788 29414 15814 29418
rect 16386 29414 16412 29440
rect 15696 29333 15722 29338
rect 15696 29316 15700 29333
rect 15700 29316 15717 29333
rect 15717 29316 15722 29333
rect 15696 29312 15722 29316
rect 15788 29312 15814 29338
rect 7048 29299 7074 29304
rect 7048 29282 7050 29299
rect 7050 29282 7074 29299
rect 7048 29278 7074 29282
rect 6956 29265 6982 29270
rect 6956 29248 6977 29265
rect 6977 29248 6982 29265
rect 10268 29278 10294 29304
rect 12108 29278 12134 29304
rect 6956 29244 6982 29248
rect 8704 29244 8730 29270
rect 8796 29244 8822 29270
rect 9026 29244 9052 29270
rect 10314 29244 10340 29270
rect 13810 29244 13836 29270
rect 14316 29244 14342 29270
rect 6726 29210 6752 29236
rect 13120 29210 13146 29236
rect 15190 29278 15216 29304
rect 13948 29176 13974 29202
rect 15788 29244 15814 29270
rect 16294 29244 16320 29270
rect 15006 29231 15032 29236
rect 15006 29214 15010 29231
rect 15010 29214 15027 29231
rect 15027 29214 15032 29231
rect 15006 29210 15032 29214
rect 15926 29231 15952 29236
rect 8060 29142 8086 29168
rect 8934 29163 8960 29168
rect 8934 29146 8938 29163
rect 8938 29146 8955 29163
rect 8955 29146 8960 29163
rect 8934 29142 8960 29146
rect 10544 29142 10570 29168
rect 11648 29142 11674 29168
rect 13902 29142 13928 29168
rect 15006 29142 15032 29168
rect 15926 29214 15930 29231
rect 15930 29214 15947 29231
rect 15947 29214 15952 29231
rect 15926 29210 15952 29214
rect 15880 29142 15906 29168
rect 6956 29040 6982 29066
rect 10360 29061 10386 29066
rect 10360 29044 10364 29061
rect 10364 29044 10381 29061
rect 10381 29044 10386 29061
rect 10360 29040 10386 29044
rect 11372 29061 11398 29066
rect 11372 29044 11376 29061
rect 11376 29044 11393 29061
rect 11393 29044 11398 29061
rect 11372 29040 11398 29044
rect 11878 29061 11904 29066
rect 11878 29044 11882 29061
rect 11882 29044 11899 29061
rect 11899 29044 11904 29061
rect 11878 29040 11904 29044
rect 13810 29040 13836 29066
rect 15190 29040 15216 29066
rect 16294 29040 16320 29066
rect 8658 29006 8684 29032
rect 8888 29006 8914 29032
rect 4702 28938 4728 28964
rect 4932 28925 4958 28930
rect 4932 28908 4936 28925
rect 4936 28908 4953 28925
rect 4953 28908 4958 28925
rect 4932 28904 4958 28908
rect 5576 28904 5602 28930
rect 6818 28938 6844 28964
rect 6864 28959 6890 28964
rect 6864 28942 6868 28959
rect 6868 28942 6885 28959
rect 6885 28942 6890 28959
rect 6864 28938 6890 28942
rect 7324 28904 7350 28930
rect 5622 28870 5648 28896
rect 7462 28959 7488 28964
rect 7462 28942 7466 28959
rect 7466 28942 7483 28959
rect 7483 28942 7488 28959
rect 7462 28938 7488 28942
rect 7508 28959 7534 28964
rect 7508 28942 7512 28959
rect 7512 28942 7529 28959
rect 7529 28942 7534 28959
rect 7508 28938 7534 28942
rect 8060 28938 8086 28964
rect 8428 28959 8454 28964
rect 8428 28942 8432 28959
rect 8432 28942 8449 28959
rect 8449 28942 8454 28959
rect 8428 28938 8454 28942
rect 8152 28904 8178 28930
rect 8934 28938 8960 28964
rect 13120 29006 13146 29032
rect 15006 29006 15032 29032
rect 15696 29027 15722 29032
rect 15696 29010 15700 29027
rect 15700 29010 15717 29027
rect 15717 29010 15722 29027
rect 15696 29006 15722 29010
rect 10406 28993 10432 28998
rect 10406 28976 10410 28993
rect 10410 28976 10427 28993
rect 10427 28976 10432 28993
rect 10406 28972 10432 28976
rect 10544 28972 10570 28998
rect 9302 28904 9328 28930
rect 10498 28938 10524 28964
rect 11188 28959 11214 28964
rect 11188 28942 11192 28959
rect 11192 28942 11209 28959
rect 11209 28942 11214 28959
rect 11188 28938 11214 28942
rect 11648 28938 11674 28964
rect 11786 28959 11812 28964
rect 11786 28942 11790 28959
rect 11790 28942 11807 28959
rect 11807 28942 11812 28959
rect 11786 28938 11812 28942
rect 13902 28972 13928 28998
rect 10360 28904 10386 28930
rect 10544 28904 10570 28930
rect 14086 28959 14112 28964
rect 14086 28942 14108 28959
rect 14108 28942 14112 28959
rect 14086 28938 14112 28942
rect 15420 28972 15446 28998
rect 14316 28870 14342 28896
rect 14592 28870 14618 28896
rect 15788 28959 15814 28964
rect 15788 28942 15792 28959
rect 15792 28942 15809 28959
rect 15809 28942 15814 28959
rect 15788 28938 15814 28942
rect 15880 28938 15906 28964
rect 16202 28959 16228 28964
rect 16202 28942 16206 28959
rect 16206 28942 16223 28959
rect 16223 28942 16228 28959
rect 16202 28938 16228 28942
rect 16248 28959 16274 28964
rect 16248 28942 16252 28959
rect 16252 28942 16269 28959
rect 16269 28942 16274 28959
rect 16248 28938 16274 28942
rect 16386 28959 16412 28964
rect 16386 28942 16390 28959
rect 16390 28942 16407 28959
rect 16407 28942 16412 28959
rect 16386 28938 16412 28942
rect 17030 28959 17056 28964
rect 17030 28942 17034 28959
rect 17034 28942 17051 28959
rect 17051 28942 17056 28959
rect 17030 28938 17056 28942
rect 17076 28959 17102 28964
rect 17076 28942 17080 28959
rect 17080 28942 17097 28959
rect 17097 28942 17102 28959
rect 17076 28938 17102 28942
rect 15742 28904 15768 28930
rect 17168 28904 17194 28930
rect 17674 28904 17700 28930
rect 17214 28891 17240 28896
rect 17214 28874 17218 28891
rect 17218 28874 17235 28891
rect 17235 28874 17240 28891
rect 17214 28870 17240 28874
rect 5530 28768 5556 28794
rect 6818 28768 6844 28794
rect 6956 28768 6982 28794
rect 8382 28768 8408 28794
rect 8428 28768 8454 28794
rect 16202 28768 16228 28794
rect 17030 28768 17056 28794
rect 18088 28768 18114 28794
rect 5990 28734 6016 28760
rect 6680 28734 6706 28760
rect 7508 28734 7534 28760
rect 5576 28700 5602 28726
rect 6588 28721 6614 28726
rect 6588 28704 6592 28721
rect 6592 28704 6609 28721
rect 6609 28704 6614 28721
rect 6588 28700 6614 28704
rect 6818 28700 6844 28726
rect 6956 28721 6982 28726
rect 6956 28704 6960 28721
rect 6960 28704 6977 28721
rect 6977 28704 6982 28721
rect 6956 28700 6982 28704
rect 7692 28700 7718 28726
rect 8658 28734 8684 28760
rect 10498 28734 10524 28760
rect 14914 28734 14940 28760
rect 20940 28768 20966 28794
rect 8152 28700 8178 28726
rect 4702 28687 4728 28692
rect 4702 28670 4706 28687
rect 4706 28670 4723 28687
rect 4723 28670 4728 28687
rect 4702 28666 4728 28670
rect 5162 28666 5188 28692
rect 8382 28700 8408 28726
rect 8796 28721 8822 28726
rect 8796 28704 8800 28721
rect 8800 28704 8817 28721
rect 8817 28704 8822 28721
rect 8796 28700 8822 28704
rect 9026 28700 9052 28726
rect 10360 28700 10386 28726
rect 8980 28666 9006 28692
rect 9348 28666 9374 28692
rect 11188 28700 11214 28726
rect 14362 28700 14388 28726
rect 15742 28700 15768 28726
rect 13258 28666 13284 28692
rect 13212 28632 13238 28658
rect 14086 28666 14112 28692
rect 15880 28721 15906 28726
rect 15880 28704 15884 28721
rect 15884 28704 15901 28721
rect 15901 28704 15906 28721
rect 15880 28700 15906 28704
rect 17398 28700 17424 28726
rect 20848 28700 20874 28726
rect 16340 28632 16366 28658
rect 16846 28632 16872 28658
rect 17214 28687 17240 28692
rect 17214 28670 17218 28687
rect 17218 28670 17235 28687
rect 17235 28670 17240 28687
rect 17214 28666 17240 28670
rect 17444 28687 17470 28692
rect 17444 28670 17448 28687
rect 17448 28670 17465 28687
rect 17465 28670 17470 28687
rect 17444 28666 17470 28670
rect 17582 28687 17608 28692
rect 17582 28670 17586 28687
rect 17586 28670 17603 28687
rect 17603 28670 17608 28687
rect 17582 28666 17608 28670
rect 20158 28687 20184 28692
rect 20158 28670 20162 28687
rect 20162 28670 20179 28687
rect 20179 28670 20184 28687
rect 20158 28666 20184 28670
rect 20296 28687 20322 28692
rect 20296 28670 20300 28687
rect 20300 28670 20317 28687
rect 20317 28670 20322 28687
rect 20296 28666 20322 28670
rect 8290 28619 8316 28624
rect 8290 28602 8294 28619
rect 8294 28602 8311 28619
rect 8311 28602 8316 28619
rect 8290 28598 8316 28602
rect 10360 28619 10386 28624
rect 10360 28602 10364 28619
rect 10364 28602 10381 28619
rect 10381 28602 10386 28619
rect 10360 28598 10386 28602
rect 13304 28598 13330 28624
rect 17260 28598 17286 28624
rect 17674 28598 17700 28624
rect 5162 28517 5188 28522
rect 5162 28500 5166 28517
rect 5166 28500 5183 28517
rect 5183 28500 5188 28517
rect 5162 28496 5188 28500
rect 5484 28449 5510 28454
rect 5484 28432 5488 28449
rect 5488 28432 5505 28449
rect 5505 28432 5510 28449
rect 6864 28483 6890 28488
rect 6864 28466 6868 28483
rect 6868 28466 6885 28483
rect 6885 28466 6890 28483
rect 6864 28462 6890 28466
rect 5484 28428 5510 28432
rect 5530 28394 5556 28420
rect 6680 28415 6706 28420
rect 6680 28398 6684 28415
rect 6684 28398 6701 28415
rect 6701 28398 6706 28415
rect 6680 28394 6706 28398
rect 6772 28415 6798 28420
rect 6772 28398 6776 28415
rect 6776 28398 6793 28415
rect 6793 28398 6798 28415
rect 6772 28394 6798 28398
rect 10222 28394 10248 28420
rect 8290 28360 8316 28386
rect 8704 28360 8730 28386
rect 10130 28360 10156 28386
rect 5530 28326 5556 28352
rect 9118 28326 9144 28352
rect 10866 28347 10892 28352
rect 10866 28330 10870 28347
rect 10870 28330 10887 28347
rect 10887 28330 10892 28347
rect 10866 28326 10892 28330
rect 14914 28394 14940 28420
rect 15466 28428 15492 28454
rect 17168 28462 17194 28488
rect 15742 28428 15768 28454
rect 15834 28394 15860 28420
rect 15972 28449 15998 28454
rect 15972 28432 15976 28449
rect 15976 28432 15993 28449
rect 15993 28432 15998 28449
rect 15972 28428 15998 28432
rect 17030 28428 17056 28454
rect 13074 28381 13100 28386
rect 13074 28364 13078 28381
rect 13078 28364 13095 28381
rect 13095 28364 13100 28381
rect 13074 28360 13100 28364
rect 13212 28360 13238 28386
rect 13120 28326 13146 28352
rect 14500 28360 14526 28386
rect 16708 28415 16734 28420
rect 16708 28398 16728 28415
rect 16728 28398 16734 28415
rect 16708 28394 16734 28398
rect 17260 28394 17286 28420
rect 20296 28517 20322 28522
rect 20296 28500 20300 28517
rect 20300 28500 20317 28517
rect 20317 28500 20322 28517
rect 20296 28496 20322 28500
rect 19238 28428 19264 28454
rect 15926 28326 15952 28352
rect 17444 28360 17470 28386
rect 16846 28347 16872 28352
rect 16846 28330 16850 28347
rect 16850 28330 16867 28347
rect 16867 28330 16872 28347
rect 18502 28360 18528 28386
rect 16846 28326 16872 28330
rect 17904 28347 17930 28352
rect 17904 28330 17908 28347
rect 17908 28330 17925 28347
rect 17925 28330 17930 28347
rect 17904 28326 17930 28330
rect 19376 28394 19402 28420
rect 20618 28428 20644 28454
rect 20894 28394 20920 28420
rect 20526 28347 20552 28352
rect 20526 28330 20530 28347
rect 20530 28330 20547 28347
rect 20547 28330 20552 28347
rect 20526 28326 20552 28330
rect 4932 28224 4958 28250
rect 5622 28224 5648 28250
rect 8980 28245 9006 28250
rect 8980 28228 8984 28245
rect 8984 28228 9001 28245
rect 9001 28228 9006 28245
rect 8980 28224 9006 28228
rect 10544 28245 10570 28250
rect 10544 28228 10548 28245
rect 10548 28228 10565 28245
rect 10565 28228 10570 28245
rect 10544 28224 10570 28228
rect 11188 28224 11214 28250
rect 13074 28224 13100 28250
rect 14500 28224 14526 28250
rect 15282 28224 15308 28250
rect 17306 28224 17332 28250
rect 17582 28224 17608 28250
rect 19376 28245 19402 28250
rect 19376 28228 19380 28245
rect 19380 28228 19397 28245
rect 19397 28228 19402 28245
rect 19376 28224 19402 28228
rect 21078 28245 21104 28250
rect 21078 28228 21082 28245
rect 21082 28228 21099 28245
rect 21099 28228 21104 28245
rect 21078 28224 21104 28228
rect 9302 28190 9328 28216
rect 5576 28156 5602 28182
rect 8750 28156 8776 28182
rect 5484 28143 5510 28148
rect 5484 28126 5488 28143
rect 5488 28126 5505 28143
rect 5505 28126 5510 28143
rect 5484 28122 5510 28126
rect 8934 28177 8960 28182
rect 8934 28160 8938 28177
rect 8938 28160 8955 28177
rect 8955 28160 8960 28177
rect 8934 28156 8960 28160
rect 9118 28156 9144 28182
rect 10176 28156 10202 28182
rect 10360 28156 10386 28182
rect 10498 28177 10524 28182
rect 10498 28160 10510 28177
rect 10510 28160 10524 28177
rect 11786 28190 11812 28216
rect 12246 28190 12272 28216
rect 10498 28156 10524 28160
rect 11004 28156 11030 28182
rect 12384 28156 12410 28182
rect 10866 28122 10892 28148
rect 11694 28122 11720 28148
rect 13304 28177 13330 28182
rect 13304 28160 13308 28177
rect 13308 28160 13325 28177
rect 13325 28160 13330 28177
rect 13304 28156 13330 28160
rect 14316 28177 14342 28182
rect 14316 28160 14320 28177
rect 14320 28160 14337 28177
rect 14337 28160 14342 28177
rect 14316 28156 14342 28160
rect 14362 28177 14388 28182
rect 14362 28160 14367 28177
rect 14367 28160 14384 28177
rect 14384 28160 14388 28177
rect 14362 28156 14388 28160
rect 14454 28177 14480 28182
rect 14454 28160 14458 28177
rect 14458 28160 14475 28177
rect 14475 28160 14480 28177
rect 14454 28156 14480 28160
rect 14500 28177 14526 28182
rect 14500 28160 14504 28177
rect 14504 28160 14521 28177
rect 14521 28160 14526 28177
rect 14500 28156 14526 28160
rect 14546 28177 14572 28182
rect 14546 28160 14553 28177
rect 14553 28160 14570 28177
rect 14570 28160 14572 28177
rect 14546 28156 14572 28160
rect 15466 28177 15492 28182
rect 15466 28160 15470 28177
rect 15470 28160 15487 28177
rect 15487 28160 15492 28177
rect 15466 28156 15492 28160
rect 15972 28190 15998 28216
rect 17398 28190 17424 28216
rect 20710 28190 20736 28216
rect 20848 28190 20874 28216
rect 15834 28177 15860 28182
rect 15834 28160 15838 28177
rect 15838 28160 15855 28177
rect 15855 28160 15860 28177
rect 15834 28156 15860 28160
rect 16708 28156 16734 28182
rect 17076 28177 17102 28182
rect 17076 28160 17080 28177
rect 17080 28160 17097 28177
rect 17097 28160 17102 28177
rect 17076 28156 17102 28160
rect 17168 28156 17194 28182
rect 17260 28156 17286 28182
rect 18088 28177 18114 28182
rect 18088 28160 18092 28177
rect 18092 28160 18109 28177
rect 18109 28160 18114 28177
rect 18088 28156 18114 28160
rect 14132 28122 14158 28148
rect 10130 28109 10156 28114
rect 10130 28092 10134 28109
rect 10134 28092 10151 28109
rect 10151 28092 10156 28109
rect 10130 28088 10156 28092
rect 17444 28088 17470 28114
rect 17812 28143 17838 28148
rect 17812 28126 17816 28143
rect 17816 28126 17833 28143
rect 17833 28126 17838 28143
rect 17812 28122 17838 28126
rect 17904 28122 17930 28148
rect 19008 28156 19034 28182
rect 18686 28143 18712 28148
rect 18686 28126 18690 28143
rect 18690 28126 18707 28143
rect 18707 28126 18712 28143
rect 18686 28122 18712 28126
rect 20158 28122 20184 28148
rect 20342 28143 20368 28148
rect 20342 28126 20346 28143
rect 20346 28126 20363 28143
rect 20363 28126 20368 28143
rect 20342 28122 20368 28126
rect 8658 28054 8684 28080
rect 10498 28054 10524 28080
rect 18088 28088 18114 28114
rect 19238 28054 19264 28080
rect 10176 27952 10202 27978
rect 17812 27952 17838 27978
rect 20342 27973 20368 27978
rect 20342 27956 20346 27973
rect 20346 27956 20363 27973
rect 20363 27956 20368 27973
rect 20342 27952 20368 27956
rect 14454 27918 14480 27944
rect 17214 27884 17240 27910
rect 17444 27905 17470 27910
rect 17444 27888 17448 27905
rect 17448 27888 17465 27905
rect 17465 27888 17470 27905
rect 17444 27884 17470 27888
rect 20618 27905 20644 27910
rect 20618 27888 20622 27905
rect 20622 27888 20639 27905
rect 20639 27888 20644 27905
rect 20618 27884 20644 27888
rect 10406 27871 10432 27876
rect 10406 27854 10410 27871
rect 10410 27854 10427 27871
rect 10427 27854 10432 27871
rect 10406 27850 10432 27854
rect 10498 27871 10524 27876
rect 10498 27854 10502 27871
rect 10502 27854 10519 27871
rect 10519 27854 10524 27871
rect 10498 27850 10524 27854
rect 11648 27850 11674 27876
rect 11786 27850 11812 27876
rect 11602 27782 11628 27808
rect 12108 27850 12134 27876
rect 12384 27871 12410 27876
rect 12384 27854 12388 27871
rect 12388 27854 12405 27871
rect 12405 27854 12410 27871
rect 12384 27850 12410 27854
rect 14500 27850 14526 27876
rect 15282 27850 15308 27876
rect 17674 27871 17700 27876
rect 17674 27854 17678 27871
rect 17678 27854 17695 27871
rect 17695 27854 17700 27871
rect 17674 27850 17700 27854
rect 18088 27850 18114 27876
rect 18686 27871 18712 27876
rect 18686 27854 18690 27871
rect 18690 27854 18707 27871
rect 18707 27854 18712 27871
rect 18686 27850 18712 27854
rect 19100 27850 19126 27876
rect 18732 27816 18758 27842
rect 17444 27782 17470 27808
rect 17904 27782 17930 27808
rect 19008 27782 19034 27808
rect 21078 27850 21104 27876
rect 19468 27782 19494 27808
rect 20572 27803 20598 27808
rect 20572 27786 20576 27803
rect 20576 27786 20593 27803
rect 20593 27786 20598 27803
rect 20572 27782 20598 27786
rect 6772 27701 6798 27706
rect 6772 27684 6776 27701
rect 6776 27684 6793 27701
rect 6793 27684 6798 27701
rect 6772 27680 6798 27684
rect 12108 27680 12134 27706
rect 4794 27646 4820 27672
rect 5070 27612 5096 27638
rect 6956 27646 6982 27672
rect 7370 27667 7396 27672
rect 7370 27650 7374 27667
rect 7374 27650 7391 27667
rect 7391 27650 7396 27667
rect 7370 27646 7396 27650
rect 8658 27646 8684 27672
rect 6680 27612 6706 27638
rect 7186 27612 7212 27638
rect 4518 27599 4544 27604
rect 4518 27582 4522 27599
rect 4522 27582 4539 27599
rect 4539 27582 4544 27599
rect 4518 27578 4544 27582
rect 5530 27578 5556 27604
rect 6956 27578 6982 27604
rect 7600 27578 7626 27604
rect 10268 27633 10294 27638
rect 10268 27616 10272 27633
rect 10272 27616 10289 27633
rect 10289 27616 10294 27633
rect 10268 27612 10294 27616
rect 10544 27646 10570 27672
rect 11648 27667 11674 27672
rect 11648 27650 11652 27667
rect 11652 27650 11669 27667
rect 11669 27650 11674 27667
rect 11648 27646 11674 27650
rect 14546 27646 14572 27672
rect 11004 27612 11030 27638
rect 11694 27633 11720 27638
rect 11694 27616 11698 27633
rect 11698 27616 11715 27633
rect 11715 27616 11720 27633
rect 11694 27612 11720 27616
rect 11924 27612 11950 27638
rect 12108 27633 12134 27638
rect 12108 27616 12112 27633
rect 12112 27616 12129 27633
rect 12129 27616 12134 27633
rect 12108 27612 12134 27616
rect 12246 27633 12272 27638
rect 12246 27616 12250 27633
rect 12250 27616 12267 27633
rect 12267 27616 12272 27633
rect 12246 27612 12272 27616
rect 13350 27633 13376 27638
rect 13350 27616 13354 27633
rect 13354 27616 13371 27633
rect 13371 27616 13376 27633
rect 13350 27612 13376 27616
rect 13396 27612 13422 27638
rect 13580 27612 13606 27638
rect 15880 27646 15906 27672
rect 17674 27646 17700 27672
rect 15144 27633 15170 27638
rect 15144 27616 15148 27633
rect 15148 27616 15165 27633
rect 15165 27616 15170 27633
rect 15144 27612 15170 27616
rect 15282 27633 15308 27638
rect 15282 27616 15286 27633
rect 15286 27616 15303 27633
rect 15303 27616 15308 27633
rect 15282 27612 15308 27616
rect 15742 27612 15768 27638
rect 17996 27633 18022 27638
rect 17996 27616 18000 27633
rect 18000 27616 18017 27633
rect 18017 27616 18022 27633
rect 17996 27612 18022 27616
rect 19238 27646 19264 27672
rect 18456 27633 18482 27638
rect 18456 27616 18460 27633
rect 18460 27616 18477 27633
rect 18477 27616 18482 27633
rect 18456 27612 18482 27616
rect 19008 27633 19034 27638
rect 19008 27616 19012 27633
rect 19012 27616 19029 27633
rect 19029 27616 19034 27633
rect 19008 27612 19034 27616
rect 7692 27578 7718 27604
rect 12338 27599 12364 27604
rect 12338 27582 12342 27599
rect 12342 27582 12359 27599
rect 12359 27582 12364 27599
rect 12338 27578 12364 27582
rect 7738 27544 7764 27570
rect 10406 27544 10432 27570
rect 10636 27544 10662 27570
rect 13304 27544 13330 27570
rect 15466 27599 15492 27604
rect 15466 27582 15470 27599
rect 15470 27582 15487 27599
rect 15487 27582 15492 27599
rect 15466 27578 15492 27582
rect 18088 27544 18114 27570
rect 18364 27544 18390 27570
rect 6358 27510 6384 27536
rect 7646 27510 7672 27536
rect 13258 27510 13284 27536
rect 18778 27544 18804 27570
rect 19376 27510 19402 27536
rect 4518 27306 4544 27332
rect 4702 27306 4728 27332
rect 6726 27408 6752 27434
rect 18732 27429 18758 27434
rect 18732 27412 18736 27429
rect 18736 27412 18753 27429
rect 18753 27412 18758 27429
rect 18732 27408 18758 27412
rect 6956 27374 6982 27400
rect 8750 27374 8776 27400
rect 14960 27395 14986 27400
rect 14960 27378 14964 27395
rect 14964 27378 14981 27395
rect 14981 27378 14986 27395
rect 14960 27374 14986 27378
rect 19468 27408 19494 27434
rect 20572 27408 20598 27434
rect 6266 27340 6292 27366
rect 7370 27340 7396 27366
rect 7646 27361 7672 27366
rect 7646 27344 7650 27361
rect 7650 27344 7667 27361
rect 7667 27344 7672 27361
rect 7646 27340 7672 27344
rect 6036 27306 6062 27332
rect 7508 27327 7534 27332
rect 7508 27310 7512 27327
rect 7512 27310 7529 27327
rect 7529 27310 7534 27327
rect 7508 27306 7534 27310
rect 7600 27327 7626 27332
rect 7600 27310 7604 27327
rect 7604 27310 7621 27327
rect 7621 27310 7626 27327
rect 7600 27306 7626 27310
rect 5622 27272 5648 27298
rect 8658 27327 8684 27332
rect 8658 27310 8662 27327
rect 8662 27310 8679 27327
rect 8679 27310 8684 27327
rect 8658 27306 8684 27310
rect 10268 27340 10294 27366
rect 9348 27327 9374 27332
rect 9348 27310 9352 27327
rect 9352 27310 9369 27327
rect 9369 27310 9374 27327
rect 9348 27306 9374 27310
rect 9716 27327 9742 27332
rect 9716 27310 9720 27327
rect 9720 27310 9737 27327
rect 9737 27310 9742 27327
rect 9716 27306 9742 27310
rect 13120 27327 13146 27332
rect 13120 27310 13124 27327
rect 13124 27310 13141 27327
rect 13141 27310 13146 27327
rect 13120 27306 13146 27310
rect 13258 27327 13284 27332
rect 13258 27310 13275 27327
rect 13275 27310 13284 27327
rect 13258 27306 13284 27310
rect 16432 27306 16458 27332
rect 8750 27293 8776 27298
rect 8750 27276 8754 27293
rect 8754 27276 8771 27293
rect 8771 27276 8776 27293
rect 8750 27272 8776 27276
rect 14592 27272 14618 27298
rect 17168 27306 17194 27332
rect 18778 27361 18804 27366
rect 18778 27344 18782 27361
rect 18782 27344 18799 27361
rect 18799 27344 18804 27361
rect 18778 27340 18804 27344
rect 6772 27238 6798 27264
rect 7048 27238 7074 27264
rect 7416 27259 7442 27264
rect 7416 27242 7420 27259
rect 7420 27242 7437 27259
rect 7437 27242 7442 27259
rect 7416 27238 7442 27242
rect 8152 27238 8178 27264
rect 13258 27238 13284 27264
rect 13396 27238 13422 27264
rect 15052 27259 15078 27264
rect 15052 27242 15056 27259
rect 15056 27242 15073 27259
rect 15073 27242 15078 27259
rect 15052 27238 15078 27242
rect 15098 27238 15124 27264
rect 16478 27238 16504 27264
rect 16570 27238 16596 27264
rect 19100 27306 19126 27332
rect 19422 27306 19448 27332
rect 19376 27293 19402 27298
rect 19376 27276 19378 27293
rect 19378 27276 19402 27293
rect 19376 27272 19402 27276
rect 5576 27136 5602 27162
rect 6036 27157 6062 27162
rect 6036 27140 6040 27157
rect 6040 27140 6057 27157
rect 6057 27140 6062 27157
rect 6036 27136 6062 27140
rect 6266 27157 6292 27162
rect 6266 27140 6270 27157
rect 6270 27140 6287 27157
rect 6287 27140 6292 27157
rect 6266 27136 6292 27140
rect 7738 27136 7764 27162
rect 11924 27157 11950 27162
rect 11924 27140 11928 27157
rect 11928 27140 11945 27157
rect 11945 27140 11950 27157
rect 11924 27136 11950 27140
rect 13350 27136 13376 27162
rect 15144 27136 15170 27162
rect 17996 27136 18022 27162
rect 5622 27102 5648 27128
rect 6772 27102 6798 27128
rect 8152 27123 8178 27128
rect 8152 27106 8156 27123
rect 8156 27106 8173 27123
rect 8173 27106 8178 27123
rect 8152 27102 8178 27106
rect 8198 27102 8224 27128
rect 9348 27102 9374 27128
rect 10636 27123 10662 27128
rect 10636 27106 10640 27123
rect 10640 27106 10657 27123
rect 10657 27106 10662 27123
rect 10636 27102 10662 27106
rect 10728 27123 10754 27128
rect 10728 27106 10740 27123
rect 10740 27106 10754 27123
rect 10728 27102 10754 27106
rect 4656 27089 4682 27094
rect 4656 27072 4677 27089
rect 4677 27072 4682 27089
rect 4656 27068 4682 27072
rect 4794 27068 4820 27094
rect 5254 27068 5280 27094
rect 6220 27089 6246 27094
rect 6220 27072 6224 27089
rect 6224 27072 6241 27089
rect 6241 27072 6246 27089
rect 6220 27068 6246 27072
rect 6726 27089 6752 27094
rect 6726 27072 6730 27089
rect 6730 27072 6747 27089
rect 6747 27072 6752 27089
rect 6726 27068 6752 27072
rect 7416 27068 7442 27094
rect 8750 27068 8776 27094
rect 11924 27068 11950 27094
rect 12384 27102 12410 27128
rect 4518 27055 4544 27060
rect 4518 27038 4522 27055
rect 4522 27038 4539 27055
rect 4539 27038 4544 27055
rect 4518 27034 4544 27038
rect 6358 27055 6384 27060
rect 6358 27038 6362 27055
rect 6362 27038 6379 27055
rect 6379 27038 6384 27055
rect 6358 27034 6384 27038
rect 7600 27034 7626 27060
rect 7416 26966 7442 26992
rect 8336 26987 8362 26992
rect 8336 26970 8340 26987
rect 8340 26970 8357 26987
rect 8357 26970 8362 26987
rect 8336 26966 8362 26970
rect 8658 26966 8684 26992
rect 12292 27089 12318 27094
rect 12292 27072 12296 27089
rect 12296 27072 12313 27089
rect 12313 27072 12318 27089
rect 14592 27102 14618 27128
rect 14960 27102 14986 27128
rect 15006 27102 15032 27128
rect 15466 27102 15492 27128
rect 16570 27102 16596 27128
rect 20710 27102 20736 27128
rect 21308 27102 21334 27128
rect 12292 27068 12318 27072
rect 13304 27068 13330 27094
rect 9716 27000 9742 27026
rect 9348 26987 9374 26992
rect 9348 26970 9352 26987
rect 9352 26970 9369 26987
rect 9369 26970 9374 26987
rect 9348 26966 9374 26970
rect 11602 27000 11628 27026
rect 13258 27034 13284 27060
rect 16340 27089 16366 27094
rect 16340 27072 16344 27089
rect 16344 27072 16361 27089
rect 16361 27072 16366 27089
rect 16340 27068 16366 27072
rect 16478 27089 16504 27094
rect 16478 27072 16482 27089
rect 16482 27072 16499 27089
rect 16499 27072 16504 27089
rect 16478 27068 16504 27072
rect 13718 27034 13744 27060
rect 14592 27055 14618 27060
rect 14592 27038 14596 27055
rect 14596 27038 14613 27055
rect 14613 27038 14618 27055
rect 14592 27034 14618 27038
rect 15098 27034 15124 27060
rect 17306 27034 17332 27060
rect 18226 27055 18252 27060
rect 18226 27038 18230 27055
rect 18230 27038 18247 27055
rect 18247 27038 18252 27055
rect 18226 27034 18252 27038
rect 18272 27055 18298 27060
rect 18272 27038 18276 27055
rect 18276 27038 18293 27055
rect 18293 27038 18298 27055
rect 18272 27034 18298 27038
rect 18364 27055 18390 27060
rect 18364 27038 18368 27055
rect 18368 27038 18385 27055
rect 18385 27038 18390 27055
rect 18364 27034 18390 27038
rect 20158 27034 20184 27060
rect 20296 27055 20322 27060
rect 20296 27038 20300 27055
rect 20300 27038 20317 27055
rect 20317 27038 20322 27055
rect 20296 27034 20322 27038
rect 20434 27055 20460 27060
rect 20434 27038 20438 27055
rect 20438 27038 20455 27055
rect 20455 27038 20460 27055
rect 20434 27034 20460 27038
rect 21124 27034 21150 27060
rect 13580 27000 13606 27026
rect 10820 26987 10846 26992
rect 10820 26970 10824 26987
rect 10824 26970 10841 26987
rect 10841 26970 10846 26987
rect 10820 26966 10846 26970
rect 11878 26966 11904 26992
rect 16616 26966 16642 26992
rect 18272 26864 18298 26890
rect 6910 26830 6936 26856
rect 7508 26830 7534 26856
rect 15052 26851 15078 26856
rect 15052 26834 15056 26851
rect 15056 26834 15073 26851
rect 15073 26834 15078 26851
rect 15052 26830 15078 26834
rect 7002 26796 7028 26822
rect 7692 26796 7718 26822
rect 8198 26796 8224 26822
rect 8658 26817 8684 26822
rect 8658 26800 8662 26817
rect 8662 26800 8679 26817
rect 8679 26800 8684 26817
rect 8658 26796 8684 26800
rect 13626 26796 13652 26822
rect 14592 26796 14618 26822
rect 18456 26796 18482 26822
rect 6634 26783 6660 26788
rect 6634 26766 6638 26783
rect 6638 26766 6655 26783
rect 6655 26766 6660 26783
rect 6634 26762 6660 26766
rect 6864 26762 6890 26788
rect 7002 26728 7028 26754
rect 7554 26783 7580 26788
rect 7554 26766 7558 26783
rect 7558 26766 7575 26783
rect 7575 26766 7580 26783
rect 7554 26762 7580 26766
rect 8612 26762 8638 26788
rect 10222 26762 10248 26788
rect 7278 26694 7304 26720
rect 8934 26728 8960 26754
rect 10820 26762 10846 26788
rect 11050 26728 11076 26754
rect 11878 26762 11904 26788
rect 12200 26783 12226 26788
rect 12200 26766 12204 26783
rect 12204 26766 12221 26783
rect 12221 26766 12226 26783
rect 12200 26762 12226 26766
rect 12292 26783 12318 26788
rect 12292 26766 12296 26783
rect 12296 26766 12313 26783
rect 12313 26766 12318 26783
rect 12292 26762 12318 26766
rect 11740 26728 11766 26754
rect 13120 26728 13146 26754
rect 13626 26728 13652 26754
rect 15144 26762 15170 26788
rect 16616 26783 16642 26788
rect 16616 26766 16633 26783
rect 16633 26766 16642 26783
rect 16616 26762 16642 26766
rect 17812 26783 17838 26788
rect 17812 26766 17816 26783
rect 17816 26766 17833 26783
rect 17833 26766 17838 26783
rect 17812 26762 17838 26766
rect 19100 26762 19126 26788
rect 17674 26728 17700 26754
rect 18640 26728 18666 26754
rect 19376 26749 19402 26754
rect 19376 26732 19378 26749
rect 19378 26732 19402 26749
rect 19376 26728 19402 26732
rect 8474 26694 8500 26720
rect 8566 26715 8592 26720
rect 8566 26698 8570 26715
rect 8570 26698 8587 26715
rect 8587 26698 8592 26715
rect 8566 26694 8592 26698
rect 10544 26694 10570 26720
rect 11970 26715 11996 26720
rect 11970 26698 11974 26715
rect 11974 26698 11991 26715
rect 11991 26698 11996 26715
rect 11970 26694 11996 26698
rect 12246 26715 12272 26720
rect 12246 26698 12250 26715
rect 12250 26698 12267 26715
rect 12267 26698 12272 26715
rect 12246 26694 12272 26698
rect 17168 26715 17194 26720
rect 17168 26698 17172 26715
rect 17172 26698 17189 26715
rect 17189 26698 17194 26715
rect 17168 26694 17194 26698
rect 17766 26694 17792 26720
rect 17904 26715 17930 26720
rect 17904 26698 17908 26715
rect 17908 26698 17925 26715
rect 17925 26698 17930 26715
rect 17904 26694 17930 26698
rect 20618 26694 20644 26720
rect 6220 26592 6246 26618
rect 6634 26592 6660 26618
rect 7186 26592 7212 26618
rect 7554 26592 7580 26618
rect 10728 26613 10754 26618
rect 10728 26596 10732 26613
rect 10732 26596 10749 26613
rect 10749 26596 10754 26613
rect 10728 26592 10754 26596
rect 6220 26545 6246 26550
rect 6220 26528 6224 26545
rect 6224 26528 6241 26545
rect 6241 26528 6246 26545
rect 6220 26524 6246 26528
rect 6956 26545 6982 26550
rect 6956 26528 6960 26545
rect 6960 26528 6977 26545
rect 6977 26528 6982 26545
rect 6956 26524 6982 26528
rect 7692 26558 7718 26584
rect 12246 26558 12272 26584
rect 17398 26592 17424 26618
rect 17812 26592 17838 26618
rect 20434 26592 20460 26618
rect 20618 26613 20644 26618
rect 20618 26596 20622 26613
rect 20622 26596 20639 26613
rect 20639 26596 20644 26613
rect 20618 26592 20644 26596
rect 15834 26558 15860 26584
rect 7186 26545 7212 26550
rect 7186 26528 7190 26545
rect 7190 26528 7207 26545
rect 7207 26528 7212 26545
rect 7186 26524 7212 26528
rect 7278 26545 7304 26550
rect 7278 26528 7282 26545
rect 7282 26528 7299 26545
rect 7299 26528 7304 26545
rect 7278 26524 7304 26528
rect 9256 26545 9282 26550
rect 9256 26528 9260 26545
rect 9260 26528 9277 26545
rect 9277 26528 9282 26545
rect 9256 26524 9282 26528
rect 10544 26545 10570 26550
rect 10544 26528 10548 26545
rect 10548 26528 10565 26545
rect 10565 26528 10570 26545
rect 10544 26524 10570 26528
rect 11740 26545 11766 26550
rect 11740 26528 11744 26545
rect 11744 26528 11761 26545
rect 11761 26528 11766 26545
rect 11740 26524 11766 26528
rect 13488 26545 13514 26550
rect 13488 26528 13492 26545
rect 13492 26528 13509 26545
rect 13509 26528 13514 26545
rect 13488 26524 13514 26528
rect 13534 26545 13560 26550
rect 13534 26528 13538 26545
rect 13538 26528 13555 26545
rect 13555 26528 13560 26545
rect 13534 26524 13560 26528
rect 13764 26524 13790 26550
rect 6864 26490 6890 26516
rect 9302 26511 9328 26516
rect 9302 26494 9306 26511
rect 9306 26494 9323 26511
rect 9323 26494 9328 26511
rect 9302 26490 9328 26494
rect 9348 26511 9374 26516
rect 9348 26494 9352 26511
rect 9352 26494 9369 26511
rect 9369 26494 9374 26511
rect 9348 26490 9374 26494
rect 10498 26511 10524 26516
rect 10498 26494 10502 26511
rect 10502 26494 10519 26511
rect 10519 26494 10524 26511
rect 10498 26490 10524 26494
rect 13580 26511 13606 26516
rect 13580 26494 13584 26511
rect 13584 26494 13601 26511
rect 13601 26494 13606 26511
rect 13580 26490 13606 26494
rect 14960 26490 14986 26516
rect 15926 26545 15952 26550
rect 15926 26528 15930 26545
rect 15930 26528 15947 26545
rect 15947 26528 15952 26545
rect 15926 26524 15952 26528
rect 17214 26558 17240 26584
rect 17168 26524 17194 26550
rect 18042 26524 18068 26550
rect 21124 26558 21150 26584
rect 18502 26524 18528 26550
rect 20250 26524 20276 26550
rect 21492 26524 21518 26550
rect 16340 26490 16366 26516
rect 17720 26490 17746 26516
rect 17904 26490 17930 26516
rect 20664 26511 20690 26516
rect 20664 26494 20668 26511
rect 20668 26494 20685 26511
rect 20685 26494 20690 26511
rect 20664 26490 20690 26494
rect 5852 26422 5878 26448
rect 9072 26443 9098 26448
rect 9072 26426 9076 26443
rect 9076 26426 9093 26443
rect 9093 26426 9098 26443
rect 9072 26422 9098 26426
rect 12476 26422 12502 26448
rect 13672 26443 13698 26448
rect 13672 26426 13676 26443
rect 13676 26426 13693 26443
rect 13693 26426 13698 26443
rect 13672 26422 13698 26426
rect 16202 26422 16228 26448
rect 16340 26422 16366 26448
rect 17858 26422 17884 26448
rect 19100 26456 19126 26482
rect 20296 26456 20322 26482
rect 22136 26422 22162 26448
rect 6220 26320 6246 26346
rect 7508 26320 7534 26346
rect 8566 26320 8592 26346
rect 12200 26320 12226 26346
rect 10820 26286 10846 26312
rect 16340 26341 16366 26346
rect 16340 26324 16344 26341
rect 16344 26324 16361 26341
rect 16361 26324 16366 26341
rect 16340 26320 16366 26324
rect 17858 26341 17884 26346
rect 17858 26324 17862 26341
rect 17862 26324 17879 26341
rect 17879 26324 17884 26341
rect 17858 26320 17884 26324
rect 17260 26286 17286 26312
rect 17996 26286 18022 26312
rect 8336 26252 8362 26278
rect 9302 26252 9328 26278
rect 5530 26239 5556 26244
rect 5530 26222 5534 26239
rect 5534 26222 5551 26239
rect 5551 26222 5556 26239
rect 5530 26218 5556 26222
rect 5852 26218 5878 26244
rect 8428 26239 8454 26244
rect 8428 26222 8432 26239
rect 8432 26222 8449 26239
rect 8449 26222 8454 26239
rect 8428 26218 8454 26222
rect 8474 26218 8500 26244
rect 11602 26239 11628 26244
rect 11602 26222 11606 26239
rect 11606 26222 11623 26239
rect 11623 26222 11628 26239
rect 11602 26218 11628 26222
rect 5576 26184 5602 26210
rect 6772 26184 6798 26210
rect 7508 26184 7534 26210
rect 7232 26150 7258 26176
rect 7554 26150 7580 26176
rect 8244 26184 8270 26210
rect 8704 26184 8730 26210
rect 12476 26218 12502 26244
rect 13028 26218 13054 26244
rect 13534 26252 13560 26278
rect 13626 26273 13652 26278
rect 13626 26256 13630 26273
rect 13630 26256 13647 26273
rect 13647 26256 13652 26273
rect 13626 26252 13652 26256
rect 14454 26252 14480 26278
rect 13258 26239 13284 26244
rect 13258 26222 13262 26239
rect 13262 26222 13279 26239
rect 13279 26222 13284 26239
rect 13258 26218 13284 26222
rect 13672 26218 13698 26244
rect 14132 26218 14158 26244
rect 14960 26273 14986 26278
rect 14960 26256 14964 26273
rect 14964 26256 14981 26273
rect 14981 26256 14986 26273
rect 14960 26252 14986 26256
rect 16294 26239 16320 26244
rect 16294 26222 16298 26239
rect 16298 26222 16315 26239
rect 16315 26222 16320 26239
rect 16294 26218 16320 26222
rect 18870 26252 18896 26278
rect 17306 26218 17332 26244
rect 19100 26239 19126 26244
rect 19100 26222 19104 26239
rect 19104 26222 19121 26239
rect 19121 26222 19126 26239
rect 19100 26218 19126 26222
rect 8934 26150 8960 26176
rect 13258 26150 13284 26176
rect 16202 26205 16228 26210
rect 16202 26188 16206 26205
rect 16206 26188 16223 26205
rect 16223 26188 16228 26205
rect 16202 26184 16228 26188
rect 17490 26184 17516 26210
rect 17720 26205 17746 26210
rect 17720 26188 17724 26205
rect 17724 26188 17741 26205
rect 17741 26188 17746 26205
rect 17720 26184 17746 26188
rect 17950 26205 17976 26210
rect 17950 26188 17954 26205
rect 17954 26188 17971 26205
rect 17971 26188 17976 26205
rect 17950 26184 17976 26188
rect 18640 26184 18666 26210
rect 19376 26218 19402 26244
rect 20526 26184 20552 26210
rect 14454 26150 14480 26176
rect 16432 26171 16458 26176
rect 16432 26154 16436 26171
rect 16436 26154 16453 26171
rect 16453 26154 16458 26171
rect 16432 26150 16458 26154
rect 17674 26150 17700 26176
rect 17996 26150 18022 26176
rect 6910 26069 6936 26074
rect 6910 26052 6914 26069
rect 6914 26052 6931 26069
rect 6931 26052 6936 26069
rect 6910 26048 6936 26052
rect 13764 26069 13790 26074
rect 13764 26052 13768 26069
rect 13768 26052 13785 26069
rect 13785 26052 13790 26069
rect 13764 26048 13790 26052
rect 18502 26069 18528 26074
rect 18502 26052 18506 26069
rect 18506 26052 18523 26069
rect 18523 26052 18528 26069
rect 18502 26048 18528 26052
rect 4472 26014 4498 26040
rect 7508 26035 7534 26040
rect 7508 26018 7510 26035
rect 7510 26018 7534 26035
rect 7508 26014 7534 26018
rect 9072 26014 9098 26040
rect 17950 26035 17976 26040
rect 17950 26018 17967 26035
rect 17967 26018 17976 26035
rect 17950 26014 17976 26018
rect 20250 26014 20276 26040
rect 22136 26014 22162 26040
rect 4840 25980 4866 26006
rect 7048 25980 7074 26006
rect 7554 25980 7580 26006
rect 8704 25980 8730 26006
rect 7002 25967 7028 25972
rect 7002 25950 7006 25967
rect 7006 25950 7023 25967
rect 7023 25950 7028 25967
rect 7002 25946 7028 25950
rect 5530 25912 5556 25938
rect 8428 25946 8454 25972
rect 8842 25946 8868 25972
rect 13028 25980 13054 26006
rect 14454 25980 14480 26006
rect 20480 25980 20506 26006
rect 21354 25980 21380 26006
rect 23010 25980 23036 26006
rect 13580 25946 13606 25972
rect 13120 25912 13146 25938
rect 13258 25912 13284 25938
rect 13718 25946 13744 25972
rect 18502 25946 18528 25972
rect 19100 25946 19126 25972
rect 21078 25946 21104 25972
rect 21584 25967 21610 25972
rect 21584 25950 21588 25967
rect 21588 25950 21605 25967
rect 21605 25950 21610 25967
rect 23286 26001 23312 26006
rect 23286 25984 23290 26001
rect 23290 25984 23307 26001
rect 23307 25984 23312 26001
rect 23286 25980 23312 25984
rect 23332 26001 23358 26006
rect 23332 25984 23336 26001
rect 23336 25984 23353 26001
rect 23353 25984 23358 26001
rect 23332 25980 23358 25984
rect 21584 25946 21610 25950
rect 23378 25967 23404 25972
rect 23378 25950 23382 25967
rect 23382 25950 23399 25967
rect 23399 25950 23404 25967
rect 23378 25946 23404 25950
rect 15006 25912 15032 25938
rect 4518 25878 4544 25904
rect 4702 25878 4728 25904
rect 6082 25878 6108 25904
rect 6634 25878 6660 25904
rect 8244 25878 8270 25904
rect 9256 25878 9282 25904
rect 10130 25878 10156 25904
rect 12982 25878 13008 25904
rect 22872 25878 22898 25904
rect 7048 25776 7074 25802
rect 7554 25776 7580 25802
rect 9256 25776 9282 25802
rect 16294 25776 16320 25802
rect 17490 25797 17516 25802
rect 17490 25780 17494 25797
rect 17494 25780 17511 25797
rect 17511 25780 17516 25797
rect 17490 25776 17516 25780
rect 23010 25797 23036 25802
rect 23010 25780 23014 25797
rect 23014 25780 23031 25797
rect 23031 25780 23036 25797
rect 23010 25776 23036 25780
rect 7232 25708 7258 25734
rect 4702 25674 4728 25700
rect 4794 25695 4820 25700
rect 4794 25678 4815 25695
rect 4815 25678 4820 25695
rect 4794 25674 4820 25678
rect 5208 25674 5234 25700
rect 7738 25695 7764 25700
rect 7738 25678 7742 25695
rect 7742 25678 7759 25695
rect 7759 25678 7764 25695
rect 7738 25674 7764 25678
rect 17122 25708 17148 25734
rect 23654 25708 23680 25734
rect 8520 25695 8546 25700
rect 8520 25678 8524 25695
rect 8524 25678 8541 25695
rect 8541 25678 8546 25695
rect 8520 25674 8546 25678
rect 6174 25606 6200 25632
rect 8106 25606 8132 25632
rect 8244 25606 8270 25632
rect 9118 25695 9144 25700
rect 9118 25678 9122 25695
rect 9122 25678 9139 25695
rect 9139 25678 9144 25695
rect 9118 25674 9144 25678
rect 9578 25674 9604 25700
rect 12982 25674 13008 25700
rect 13488 25674 13514 25700
rect 13534 25640 13560 25666
rect 16708 25674 16734 25700
rect 17214 25674 17240 25700
rect 20480 25674 20506 25700
rect 21538 25674 21564 25700
rect 17260 25640 17286 25666
rect 22872 25695 22898 25700
rect 22872 25678 22876 25695
rect 22876 25678 22893 25695
rect 22893 25678 22898 25695
rect 22872 25674 22898 25678
rect 23102 25695 23128 25700
rect 23102 25678 23106 25695
rect 23106 25678 23123 25695
rect 23123 25678 23128 25695
rect 23102 25674 23128 25678
rect 15926 25606 15952 25632
rect 21354 25606 21380 25632
rect 21446 25606 21472 25632
rect 21584 25606 21610 25632
rect 4886 25504 4912 25530
rect 5530 25504 5556 25530
rect 7554 25504 7580 25530
rect 8520 25504 8546 25530
rect 8658 25504 8684 25530
rect 8842 25504 8868 25530
rect 9624 25504 9650 25530
rect 18870 25525 18896 25530
rect 18870 25508 18874 25525
rect 18874 25508 18891 25525
rect 18891 25508 18896 25525
rect 18870 25504 18896 25508
rect 23654 25525 23680 25530
rect 23654 25508 23658 25525
rect 23658 25508 23675 25525
rect 23675 25508 23680 25525
rect 23654 25504 23680 25508
rect 3276 25470 3302 25496
rect 3414 25436 3440 25462
rect 6772 25470 6798 25496
rect 3644 25436 3670 25462
rect 5530 25436 5556 25462
rect 6634 25457 6660 25462
rect 6634 25440 6655 25457
rect 6655 25440 6660 25457
rect 6634 25436 6660 25440
rect 7416 25402 7442 25428
rect 8336 25402 8362 25428
rect 8934 25402 8960 25428
rect 4472 25368 4498 25394
rect 4794 25334 4820 25360
rect 8060 25368 8086 25394
rect 8152 25368 8178 25394
rect 9072 25436 9098 25462
rect 18318 25470 18344 25496
rect 10682 25436 10708 25462
rect 17904 25436 17930 25462
rect 18778 25436 18804 25462
rect 9624 25334 9650 25360
rect 18916 25402 18942 25428
rect 23332 25436 23358 25462
rect 23286 25402 23312 25428
rect 11050 25368 11076 25394
rect 23102 25368 23128 25394
rect 10774 25334 10800 25360
rect 19100 25355 19126 25360
rect 19100 25338 19104 25355
rect 19104 25338 19121 25355
rect 19121 25338 19126 25355
rect 19100 25334 19126 25338
rect 23562 25355 23588 25360
rect 23562 25338 23566 25355
rect 23566 25338 23583 25355
rect 23583 25338 23588 25355
rect 23562 25334 23588 25338
rect 3414 25232 3440 25258
rect 8152 25232 8178 25258
rect 11234 25232 11260 25258
rect 12844 25232 12870 25258
rect 17398 25253 17424 25258
rect 17398 25236 17402 25253
rect 17402 25236 17419 25253
rect 17419 25236 17424 25253
rect 17398 25232 17424 25236
rect 23102 25232 23128 25258
rect 3276 25151 3302 25156
rect 3276 25134 3297 25151
rect 3297 25134 3302 25151
rect 3276 25130 3302 25134
rect 3736 25130 3762 25156
rect 4794 25151 4820 25156
rect 4794 25134 4798 25151
rect 4798 25134 4815 25151
rect 4815 25134 4820 25151
rect 4794 25130 4820 25134
rect 5254 25130 5280 25156
rect 8290 25130 8316 25156
rect 8658 25151 8684 25156
rect 8658 25134 8662 25151
rect 8662 25134 8679 25151
rect 8679 25134 8684 25151
rect 8658 25130 8684 25134
rect 4886 25096 4912 25122
rect 8336 25096 8362 25122
rect 11004 25151 11030 25156
rect 11004 25134 11008 25151
rect 11008 25134 11025 25151
rect 11025 25134 11030 25151
rect 11004 25130 11030 25134
rect 11326 25130 11352 25156
rect 15052 25164 15078 25190
rect 17076 25164 17102 25190
rect 18364 25164 18390 25190
rect 18502 25185 18528 25190
rect 18502 25168 18506 25185
rect 18506 25168 18523 25185
rect 18523 25168 18528 25185
rect 18502 25164 18528 25168
rect 14914 25151 14940 25156
rect 14914 25134 14918 25151
rect 14918 25134 14935 25151
rect 14935 25134 14940 25151
rect 14914 25130 14940 25134
rect 15006 25130 15032 25156
rect 16156 25130 16182 25156
rect 11234 25117 11260 25122
rect 11234 25100 11236 25117
rect 11236 25100 11260 25117
rect 11234 25096 11260 25100
rect 6358 25062 6384 25088
rect 10498 25062 10524 25088
rect 12062 25062 12088 25088
rect 14500 25062 14526 25088
rect 17168 25096 17194 25122
rect 19100 25130 19126 25156
rect 20480 25130 20506 25156
rect 21676 25151 21702 25156
rect 21676 25134 21680 25151
rect 21680 25134 21697 25151
rect 21697 25134 21702 25151
rect 21676 25130 21702 25134
rect 23930 25130 23956 25156
rect 17720 25117 17746 25122
rect 17720 25100 17724 25117
rect 17724 25100 17741 25117
rect 17741 25100 17746 25117
rect 17720 25096 17746 25100
rect 18548 25096 18574 25122
rect 21906 25117 21932 25122
rect 18686 25062 18712 25088
rect 21906 25100 21908 25117
rect 21908 25100 21932 25117
rect 21906 25096 21932 25100
rect 20388 25062 20414 25088
rect 9670 24926 9696 24952
rect 10682 24926 10708 24952
rect 5806 24892 5832 24918
rect 6082 24913 6108 24918
rect 6082 24896 6097 24913
rect 6097 24896 6108 24913
rect 6082 24892 6108 24896
rect 6174 24913 6200 24918
rect 6174 24896 6191 24913
rect 6191 24896 6200 24913
rect 6174 24892 6200 24896
rect 7784 24892 7810 24918
rect 8934 24892 8960 24918
rect 11372 24892 11398 24918
rect 12798 24892 12824 24918
rect 6542 24858 6568 24884
rect 9624 24879 9650 24884
rect 9624 24862 9628 24879
rect 9628 24862 9645 24879
rect 9645 24862 9650 24879
rect 9624 24858 9650 24862
rect 11050 24858 11076 24884
rect 6496 24824 6522 24850
rect 13120 24913 13146 24918
rect 13120 24896 13124 24913
rect 13124 24896 13141 24913
rect 13141 24896 13146 24913
rect 13120 24892 13146 24896
rect 13258 24913 13284 24918
rect 13258 24896 13262 24913
rect 13262 24896 13279 24913
rect 13279 24896 13284 24913
rect 13258 24892 13284 24896
rect 13994 24892 14020 24918
rect 14776 24892 14802 24918
rect 15006 24960 15032 24986
rect 15880 24960 15906 24986
rect 18318 24960 18344 24986
rect 14914 24926 14940 24952
rect 15052 24858 15078 24884
rect 15880 24913 15906 24918
rect 15880 24896 15884 24913
rect 15884 24896 15901 24913
rect 15901 24896 15906 24913
rect 15880 24892 15906 24896
rect 17076 24913 17102 24918
rect 17076 24896 17080 24913
rect 17080 24896 17097 24913
rect 17097 24896 17102 24913
rect 17076 24892 17102 24896
rect 17260 24892 17286 24918
rect 18548 24892 18574 24918
rect 17168 24858 17194 24884
rect 18318 24879 18344 24884
rect 18318 24862 18322 24879
rect 18322 24862 18339 24879
rect 18339 24862 18344 24879
rect 18318 24858 18344 24862
rect 18456 24858 18482 24884
rect 18686 24879 18712 24884
rect 18686 24862 18690 24879
rect 18690 24862 18707 24879
rect 18707 24862 18712 24879
rect 18686 24858 18712 24862
rect 18916 24879 18942 24884
rect 18916 24862 18920 24879
rect 18920 24862 18937 24879
rect 18937 24862 18942 24879
rect 18916 24858 18942 24862
rect 20388 24879 20414 24884
rect 20388 24862 20392 24879
rect 20392 24862 20409 24879
rect 20409 24862 20414 24879
rect 20388 24858 20414 24862
rect 6404 24790 6430 24816
rect 10636 24790 10662 24816
rect 11326 24790 11352 24816
rect 13810 24824 13836 24850
rect 18778 24824 18804 24850
rect 21400 24913 21426 24918
rect 21400 24896 21404 24913
rect 21404 24896 21421 24913
rect 21421 24896 21426 24913
rect 21400 24892 21426 24896
rect 21538 24858 21564 24884
rect 12430 24790 12456 24816
rect 14408 24790 14434 24816
rect 14868 24811 14894 24816
rect 14868 24794 14872 24811
rect 14872 24794 14889 24811
rect 14889 24794 14894 24811
rect 14868 24790 14894 24794
rect 16018 24811 16044 24816
rect 16018 24794 16022 24811
rect 16022 24794 16039 24811
rect 16039 24794 16044 24811
rect 16018 24790 16044 24794
rect 17122 24811 17148 24816
rect 17122 24794 17126 24811
rect 17126 24794 17143 24811
rect 17143 24794 17148 24811
rect 17122 24790 17148 24794
rect 20342 24790 20368 24816
rect 5806 24688 5832 24714
rect 6542 24688 6568 24714
rect 10728 24654 10754 24680
rect 10774 24654 10800 24680
rect 6956 24620 6982 24646
rect 5162 24586 5188 24612
rect 5530 24607 5556 24612
rect 5530 24590 5534 24607
rect 5534 24590 5551 24607
rect 5551 24590 5556 24607
rect 5530 24586 5556 24590
rect 5668 24607 5694 24612
rect 5668 24590 5689 24607
rect 5689 24590 5694 24607
rect 5668 24586 5694 24590
rect 6220 24586 6246 24612
rect 7922 24607 7948 24612
rect 7922 24590 7929 24607
rect 7929 24590 7946 24607
rect 7946 24590 7948 24607
rect 7922 24586 7948 24590
rect 8198 24607 8224 24612
rect 8198 24590 8202 24607
rect 8202 24590 8219 24607
rect 8219 24590 8224 24607
rect 8198 24586 8224 24590
rect 8244 24586 8270 24612
rect 9210 24586 9236 24612
rect 10498 24607 10524 24612
rect 10498 24590 10502 24607
rect 10502 24590 10519 24607
rect 10519 24590 10524 24607
rect 10498 24586 10524 24590
rect 10544 24607 10570 24612
rect 10544 24590 10559 24607
rect 10559 24590 10570 24607
rect 10544 24586 10570 24590
rect 10636 24605 10662 24612
rect 10636 24588 10653 24605
rect 10653 24588 10662 24605
rect 12338 24688 12364 24714
rect 18226 24688 18252 24714
rect 23332 24688 23358 24714
rect 23654 24688 23680 24714
rect 12384 24620 12410 24646
rect 14776 24641 14802 24646
rect 14776 24624 14780 24641
rect 14780 24624 14797 24641
rect 14797 24624 14802 24641
rect 14776 24620 14802 24624
rect 14914 24620 14940 24646
rect 15052 24641 15078 24646
rect 15052 24624 15056 24641
rect 15056 24624 15073 24641
rect 15073 24624 15078 24641
rect 15052 24620 15078 24624
rect 10636 24586 10662 24588
rect 11050 24586 11076 24612
rect 11372 24586 11398 24612
rect 12982 24586 13008 24612
rect 7738 24573 7764 24578
rect 7738 24556 7742 24573
rect 7742 24556 7759 24573
rect 7759 24556 7764 24573
rect 7738 24552 7764 24556
rect 7876 24573 7902 24578
rect 7876 24556 7880 24573
rect 7880 24556 7897 24573
rect 7897 24556 7902 24573
rect 7876 24552 7902 24556
rect 11326 24573 11352 24578
rect 11326 24556 11328 24573
rect 11328 24556 11352 24573
rect 11326 24552 11352 24556
rect 13810 24586 13836 24612
rect 13994 24586 14020 24612
rect 14500 24586 14526 24612
rect 14822 24586 14848 24612
rect 14868 24586 14894 24612
rect 16708 24607 16734 24612
rect 16708 24590 16712 24607
rect 16712 24590 16729 24607
rect 16729 24590 16734 24607
rect 16708 24586 16734 24590
rect 17260 24620 17286 24646
rect 18594 24641 18620 24646
rect 18594 24624 18598 24641
rect 18598 24624 18615 24641
rect 18615 24624 18620 24641
rect 18594 24620 18620 24624
rect 19422 24620 19448 24646
rect 17076 24607 17102 24612
rect 17076 24590 17080 24607
rect 17080 24590 17097 24607
rect 17097 24590 17102 24607
rect 17076 24586 17102 24590
rect 17904 24586 17930 24612
rect 18548 24607 18574 24612
rect 18548 24590 18552 24607
rect 18552 24590 18569 24607
rect 18569 24590 18574 24607
rect 18548 24586 18574 24590
rect 19560 24607 19586 24612
rect 19560 24590 19564 24607
rect 19564 24590 19581 24607
rect 19581 24590 19586 24607
rect 19560 24586 19586 24590
rect 20250 24586 20276 24612
rect 21906 24620 21932 24646
rect 21676 24586 21702 24612
rect 15650 24552 15676 24578
rect 8060 24518 8086 24544
rect 8244 24518 8270 24544
rect 9302 24518 9328 24544
rect 10682 24518 10708 24544
rect 12154 24518 12180 24544
rect 12798 24518 12824 24544
rect 13672 24539 13698 24544
rect 13672 24522 13676 24539
rect 13676 24522 13693 24539
rect 13693 24522 13698 24539
rect 13672 24518 13698 24522
rect 15052 24518 15078 24544
rect 19606 24552 19632 24578
rect 21998 24552 22024 24578
rect 23930 24586 23956 24612
rect 24068 24573 24094 24578
rect 24068 24556 24072 24573
rect 24072 24556 24089 24573
rect 24089 24556 24094 24573
rect 24068 24552 24094 24556
rect 20388 24518 20414 24544
rect 7738 24416 7764 24442
rect 8014 24416 8040 24442
rect 10728 24416 10754 24442
rect 12108 24416 12134 24442
rect 13994 24416 14020 24442
rect 14178 24416 14204 24442
rect 16156 24416 16182 24442
rect 17766 24437 17792 24442
rect 17766 24420 17770 24437
rect 17770 24420 17787 24437
rect 17787 24420 17792 24437
rect 17766 24416 17792 24420
rect 8060 24382 8086 24408
rect 9302 24403 9328 24408
rect 9302 24386 9306 24403
rect 9306 24386 9323 24403
rect 9323 24386 9328 24403
rect 9302 24382 9328 24386
rect 3276 24348 3302 24374
rect 3506 24348 3532 24374
rect 5852 24348 5878 24374
rect 7048 24369 7074 24374
rect 7048 24352 7069 24369
rect 7069 24352 7074 24369
rect 7048 24348 7074 24352
rect 7554 24348 7580 24374
rect 9164 24369 9190 24374
rect 9164 24352 9168 24369
rect 9168 24352 9185 24369
rect 9185 24352 9190 24369
rect 9164 24348 9190 24352
rect 9256 24369 9282 24374
rect 9256 24352 9260 24369
rect 9260 24352 9277 24369
rect 9277 24352 9282 24369
rect 9256 24348 9282 24352
rect 9348 24369 9374 24374
rect 9348 24352 9355 24369
rect 9355 24352 9372 24369
rect 9372 24352 9374 24369
rect 9348 24348 9374 24352
rect 10544 24348 10570 24374
rect 12016 24369 12042 24374
rect 12016 24352 12020 24369
rect 12020 24352 12037 24369
rect 12037 24352 12042 24369
rect 12016 24348 12042 24352
rect 12062 24369 12088 24374
rect 12062 24352 12077 24369
rect 12077 24352 12088 24369
rect 12062 24348 12088 24352
rect 12154 24369 12180 24374
rect 12154 24352 12171 24369
rect 12171 24352 12180 24369
rect 12430 24382 12456 24408
rect 14914 24382 14940 24408
rect 16018 24382 16044 24408
rect 12338 24369 12364 24374
rect 12154 24348 12180 24352
rect 12338 24352 12349 24369
rect 12349 24352 12364 24369
rect 12338 24348 12364 24352
rect 15144 24348 15170 24374
rect 3414 24314 3440 24340
rect 6910 24335 6936 24340
rect 6910 24318 6914 24335
rect 6914 24318 6931 24335
rect 6931 24318 6936 24335
rect 6910 24314 6936 24318
rect 9440 24314 9466 24340
rect 13810 24314 13836 24340
rect 13994 24314 14020 24340
rect 14454 24314 14480 24340
rect 16156 24369 16182 24374
rect 16156 24352 16160 24369
rect 16160 24352 16177 24369
rect 16177 24352 16182 24369
rect 16156 24348 16182 24352
rect 17720 24348 17746 24374
rect 19606 24348 19632 24374
rect 17536 24335 17562 24340
rect 17536 24318 17540 24335
rect 17540 24318 17557 24335
rect 17557 24318 17562 24335
rect 17536 24314 17562 24318
rect 20388 24335 20414 24340
rect 20388 24318 20392 24335
rect 20392 24318 20409 24335
rect 20409 24318 20414 24335
rect 20388 24314 20414 24318
rect 21078 24416 21104 24442
rect 23562 24416 23588 24442
rect 22826 24382 22852 24408
rect 20986 24369 21012 24374
rect 20986 24352 20990 24369
rect 20990 24352 21007 24369
rect 21007 24352 21012 24369
rect 20986 24348 21012 24352
rect 12384 24280 12410 24306
rect 16340 24301 16366 24306
rect 16340 24284 16344 24301
rect 16344 24284 16361 24301
rect 16361 24284 16366 24301
rect 16340 24280 16366 24284
rect 5024 24246 5050 24272
rect 6496 24246 6522 24272
rect 9348 24246 9374 24272
rect 9624 24246 9650 24272
rect 12154 24246 12180 24272
rect 22090 24348 22116 24374
rect 22964 24369 22990 24374
rect 22964 24352 22968 24369
rect 22968 24352 22985 24369
rect 22985 24352 22990 24369
rect 22964 24348 22990 24352
rect 23240 24348 23266 24374
rect 23378 24369 23404 24374
rect 23378 24352 23382 24369
rect 23382 24352 23399 24369
rect 23399 24352 23404 24369
rect 23378 24348 23404 24352
rect 23470 24403 23496 24408
rect 23470 24386 23484 24403
rect 23484 24386 23496 24403
rect 23470 24382 23496 24386
rect 24114 24382 24140 24408
rect 23746 24348 23772 24374
rect 21170 24335 21196 24340
rect 21170 24318 21174 24335
rect 21174 24318 21191 24335
rect 21191 24318 21196 24335
rect 21170 24314 21196 24318
rect 22918 24335 22944 24340
rect 22918 24318 22922 24335
rect 22922 24318 22939 24335
rect 22939 24318 22944 24335
rect 22918 24314 22944 24318
rect 24068 24369 24094 24374
rect 24068 24352 24072 24369
rect 24072 24352 24089 24369
rect 24089 24352 24094 24369
rect 24068 24348 24094 24352
rect 24114 24314 24140 24340
rect 23286 24280 23312 24306
rect 24620 24280 24646 24306
rect 23930 24267 23956 24272
rect 23930 24250 23934 24267
rect 23934 24250 23951 24267
rect 23951 24250 23956 24267
rect 23930 24246 23956 24250
rect 3414 24144 3440 24170
rect 5070 24110 5096 24136
rect 5530 24110 5556 24136
rect 5668 24110 5694 24136
rect 7048 24110 7074 24136
rect 6910 24076 6936 24102
rect 8198 24144 8224 24170
rect 9164 24144 9190 24170
rect 9210 24144 9236 24170
rect 13212 24144 13238 24170
rect 13672 24144 13698 24170
rect 22918 24144 22944 24170
rect 9026 24110 9052 24136
rect 16294 24076 16320 24102
rect 17122 24076 17148 24102
rect 18456 24131 18482 24136
rect 18456 24114 18460 24131
rect 18460 24114 18477 24131
rect 18477 24114 18482 24131
rect 18456 24110 18482 24114
rect 20986 24110 21012 24136
rect 24436 24110 24462 24136
rect 18640 24076 18666 24102
rect 20434 24097 20460 24102
rect 20434 24080 20438 24097
rect 20438 24080 20455 24097
rect 20455 24080 20460 24097
rect 20434 24076 20460 24080
rect 21676 24076 21702 24102
rect 24252 24097 24278 24102
rect 24252 24080 24256 24097
rect 24256 24080 24273 24097
rect 24273 24080 24278 24097
rect 24252 24076 24278 24080
rect 3460 24042 3486 24068
rect 4932 24042 4958 24068
rect 8336 24042 8362 24068
rect 9164 24042 9190 24068
rect 12154 24063 12180 24068
rect 12154 24046 12158 24063
rect 12158 24046 12175 24063
rect 12175 24046 12180 24063
rect 12154 24042 12180 24046
rect 12292 24063 12318 24068
rect 12292 24046 12296 24063
rect 12296 24046 12313 24063
rect 12313 24046 12318 24063
rect 12292 24042 12318 24046
rect 12660 24042 12686 24068
rect 13994 24063 14020 24068
rect 13994 24046 13998 24063
rect 13998 24046 14015 24063
rect 14015 24046 14020 24063
rect 13994 24042 14020 24046
rect 14178 24063 14204 24068
rect 14178 24046 14182 24063
rect 14182 24046 14199 24063
rect 14199 24046 14204 24063
rect 14178 24042 14204 24046
rect 14500 24042 14526 24068
rect 14868 24042 14894 24068
rect 16340 24063 16366 24068
rect 16340 24046 16344 24063
rect 16344 24046 16361 24063
rect 16361 24046 16366 24063
rect 16340 24042 16366 24046
rect 16708 24042 16734 24068
rect 17904 24042 17930 24068
rect 18088 24042 18114 24068
rect 18594 24063 18620 24068
rect 18594 24046 18598 24063
rect 18598 24046 18615 24063
rect 18615 24046 18620 24063
rect 18594 24042 18620 24046
rect 20020 24042 20046 24068
rect 21400 24042 21426 24068
rect 23240 24042 23266 24068
rect 24114 24063 24140 24068
rect 24114 24046 24118 24063
rect 24118 24046 24135 24063
rect 24135 24046 24140 24063
rect 24114 24042 24140 24046
rect 3184 24008 3210 24034
rect 3368 24029 3394 24034
rect 3368 24012 3370 24029
rect 3370 24012 3394 24029
rect 3368 24008 3394 24012
rect 4748 23974 4774 24000
rect 6956 24008 6982 24034
rect 7554 24008 7580 24034
rect 18502 24008 18528 24034
rect 21952 24029 21978 24034
rect 21952 24012 21954 24029
rect 21954 24012 21978 24029
rect 21952 24008 21978 24012
rect 24620 24063 24646 24068
rect 24620 24046 24624 24063
rect 24624 24046 24641 24063
rect 24641 24046 24646 24063
rect 24620 24042 24646 24046
rect 24804 24008 24830 24034
rect 5576 23974 5602 24000
rect 13902 23995 13928 24000
rect 13902 23978 13906 23995
rect 13906 23978 13923 23995
rect 13923 23978 13928 23995
rect 13902 23974 13928 23978
rect 16386 23995 16412 24000
rect 16386 23978 16390 23995
rect 16390 23978 16407 23995
rect 16407 23978 16412 23995
rect 16386 23974 16412 23978
rect 17030 23974 17056 24000
rect 17996 23974 18022 24000
rect 18594 23974 18620 24000
rect 23608 23974 23634 24000
rect 24114 23974 24140 24000
rect 4840 23872 4866 23898
rect 4932 23872 4958 23898
rect 5024 23872 5050 23898
rect 17904 23872 17930 23898
rect 21584 23872 21610 23898
rect 23746 23893 23772 23898
rect 23746 23876 23750 23893
rect 23750 23876 23767 23893
rect 23767 23876 23772 23893
rect 23746 23872 23772 23876
rect 3460 23838 3486 23864
rect 3690 23859 3716 23864
rect 3690 23842 3692 23859
rect 3692 23842 3716 23859
rect 3690 23838 3716 23842
rect 4748 23825 4774 23830
rect 4748 23808 4752 23825
rect 4752 23808 4769 23825
rect 4769 23808 4774 23825
rect 4748 23804 4774 23808
rect 6358 23859 6384 23864
rect 6358 23842 6362 23859
rect 6362 23842 6379 23859
rect 6379 23842 6384 23859
rect 6358 23838 6384 23842
rect 6956 23838 6982 23864
rect 3414 23770 3440 23796
rect 4886 23736 4912 23762
rect 6450 23825 6476 23830
rect 6450 23808 6454 23825
rect 6454 23808 6471 23825
rect 6471 23808 6476 23825
rect 6450 23804 6476 23808
rect 6818 23804 6844 23830
rect 6910 23825 6936 23830
rect 6910 23808 6914 23825
rect 6914 23808 6931 23825
rect 6931 23808 6936 23825
rect 6910 23804 6936 23808
rect 7048 23804 7074 23830
rect 7324 23804 7350 23830
rect 6588 23770 6614 23796
rect 3644 23702 3670 23728
rect 5254 23702 5280 23728
rect 6036 23702 6062 23728
rect 6358 23723 6384 23728
rect 6358 23706 6362 23723
rect 6362 23706 6379 23723
rect 6379 23706 6384 23723
rect 6358 23702 6384 23706
rect 9026 23825 9052 23830
rect 9026 23808 9030 23825
rect 9030 23808 9047 23825
rect 9047 23808 9052 23825
rect 9026 23804 9052 23808
rect 9164 23825 9190 23830
rect 9164 23808 9185 23825
rect 9185 23808 9190 23825
rect 9164 23804 9190 23808
rect 11326 23804 11352 23830
rect 13120 23838 13146 23864
rect 13534 23838 13560 23864
rect 13258 23804 13284 23830
rect 7876 23770 7902 23796
rect 13304 23770 13330 23796
rect 14960 23825 14986 23830
rect 14960 23808 14964 23825
rect 14964 23808 14981 23825
rect 14981 23808 14986 23825
rect 14960 23804 14986 23808
rect 15052 23825 15078 23830
rect 15052 23808 15056 23825
rect 15056 23808 15073 23825
rect 15073 23808 15078 23825
rect 15052 23804 15078 23808
rect 18456 23859 18482 23864
rect 18456 23842 18473 23859
rect 18473 23842 18482 23859
rect 18456 23838 18482 23842
rect 21676 23838 21702 23864
rect 18364 23804 18390 23830
rect 19376 23804 19402 23830
rect 19560 23804 19586 23830
rect 21446 23825 21472 23830
rect 21446 23808 21450 23825
rect 21450 23808 21467 23825
rect 21467 23808 21472 23825
rect 21446 23804 21472 23808
rect 24252 23872 24278 23898
rect 23930 23838 23956 23864
rect 15190 23791 15216 23796
rect 15190 23774 15194 23791
rect 15194 23774 15211 23791
rect 15211 23774 15216 23791
rect 15190 23770 15216 23774
rect 17950 23791 17976 23796
rect 17950 23774 17954 23791
rect 17954 23774 17971 23791
rect 17971 23774 17976 23791
rect 17950 23770 17976 23774
rect 18088 23791 18114 23796
rect 18088 23774 18092 23791
rect 18092 23774 18109 23791
rect 18109 23774 18114 23791
rect 18088 23770 18114 23774
rect 21308 23770 21334 23796
rect 23608 23791 23634 23796
rect 23608 23774 23612 23791
rect 23612 23774 23629 23791
rect 23629 23774 23634 23791
rect 23608 23770 23634 23774
rect 24390 23804 24416 23830
rect 9670 23702 9696 23728
rect 10958 23736 10984 23762
rect 14638 23736 14664 23762
rect 10222 23702 10248 23728
rect 21492 23702 21518 23728
rect 24528 23702 24554 23728
rect 5070 23600 5096 23626
rect 5254 23600 5280 23626
rect 5576 23600 5602 23626
rect 6404 23587 6430 23592
rect 6404 23570 6408 23587
rect 6408 23570 6425 23587
rect 6425 23570 6430 23587
rect 6404 23566 6430 23570
rect 6036 23532 6062 23558
rect 3414 23498 3440 23524
rect 5162 23498 5188 23524
rect 3460 23464 3486 23490
rect 5530 23498 5556 23524
rect 6358 23498 6384 23524
rect 8152 23519 8178 23524
rect 8152 23502 8156 23519
rect 8156 23502 8173 23519
rect 8173 23502 8178 23519
rect 8152 23498 8178 23502
rect 8290 23519 8316 23524
rect 8290 23502 8311 23519
rect 8311 23502 8316 23519
rect 8290 23498 8316 23502
rect 8888 23498 8914 23524
rect 9440 23519 9466 23524
rect 9440 23502 9444 23519
rect 9444 23502 9461 23519
rect 9461 23502 9466 23519
rect 9440 23498 9466 23502
rect 9532 23519 9558 23524
rect 9532 23502 9536 23519
rect 9536 23502 9553 23519
rect 9553 23502 9558 23519
rect 9532 23498 9558 23502
rect 10222 23519 10248 23524
rect 10222 23502 10226 23519
rect 10226 23502 10243 23519
rect 10243 23502 10248 23519
rect 10222 23498 10248 23502
rect 12384 23600 12410 23626
rect 18502 23600 18528 23626
rect 20434 23600 20460 23626
rect 17904 23566 17930 23592
rect 10958 23532 10984 23558
rect 10406 23519 10432 23524
rect 10406 23502 10410 23519
rect 10410 23502 10427 23519
rect 10427 23502 10432 23519
rect 10406 23498 10432 23502
rect 11004 23519 11030 23524
rect 11004 23502 11008 23519
rect 11008 23502 11025 23519
rect 11025 23502 11030 23519
rect 11004 23498 11030 23502
rect 17076 23532 17102 23558
rect 5346 23485 5372 23490
rect 5346 23468 5348 23485
rect 5348 23468 5372 23485
rect 5346 23464 5372 23468
rect 8382 23485 8408 23490
rect 8382 23468 8384 23485
rect 8384 23468 8408 23485
rect 8382 23464 8408 23468
rect 10360 23485 10386 23490
rect 10360 23468 10364 23485
rect 10364 23468 10381 23485
rect 10381 23468 10386 23485
rect 10360 23464 10386 23468
rect 11418 23498 11444 23524
rect 12982 23519 13008 23524
rect 12982 23502 12986 23519
rect 12986 23502 13003 23519
rect 13003 23502 13008 23519
rect 12982 23498 13008 23502
rect 13258 23519 13284 23524
rect 13258 23502 13262 23519
rect 13262 23502 13279 23519
rect 13279 23502 13284 23519
rect 13258 23498 13284 23502
rect 16708 23498 16734 23524
rect 17950 23532 17976 23558
rect 18134 23532 18160 23558
rect 21216 23587 21242 23592
rect 21216 23570 21220 23587
rect 21220 23570 21237 23587
rect 21237 23570 21242 23587
rect 21216 23566 21242 23570
rect 22688 23566 22714 23592
rect 23608 23566 23634 23592
rect 18548 23532 18574 23558
rect 19376 23553 19402 23558
rect 19376 23536 19380 23553
rect 19380 23536 19397 23553
rect 19397 23536 19402 23553
rect 19376 23532 19402 23536
rect 21400 23532 21426 23558
rect 21722 23532 21748 23558
rect 17260 23464 17286 23490
rect 17812 23464 17838 23490
rect 20020 23498 20046 23524
rect 21354 23519 21380 23524
rect 21354 23502 21358 23519
rect 21358 23502 21375 23519
rect 21375 23502 21380 23519
rect 21354 23498 21380 23502
rect 21952 23498 21978 23524
rect 23424 23498 23450 23524
rect 24436 23519 24462 23524
rect 24436 23502 24453 23519
rect 24453 23502 24462 23519
rect 18594 23464 18620 23490
rect 19422 23464 19448 23490
rect 21262 23464 21288 23490
rect 22044 23485 22070 23490
rect 22044 23468 22046 23485
rect 22046 23468 22070 23485
rect 22044 23464 22070 23468
rect 24436 23498 24462 23502
rect 24390 23464 24416 23490
rect 6266 23430 6292 23456
rect 6312 23430 6338 23456
rect 8198 23430 8224 23456
rect 9394 23430 9420 23456
rect 10636 23430 10662 23456
rect 12016 23430 12042 23456
rect 12890 23430 12916 23456
rect 15236 23430 15262 23456
rect 15834 23430 15860 23456
rect 17950 23430 17976 23456
rect 21584 23430 21610 23456
rect 23378 23451 23404 23456
rect 23378 23434 23382 23451
rect 23382 23434 23399 23451
rect 23399 23434 23404 23451
rect 23378 23430 23404 23434
rect 24804 23430 24830 23456
rect 10360 23328 10386 23354
rect 10682 23349 10708 23354
rect 10682 23332 10686 23349
rect 10686 23332 10703 23349
rect 10703 23332 10708 23349
rect 10682 23328 10708 23332
rect 10728 23349 10754 23354
rect 10728 23332 10732 23349
rect 10732 23332 10749 23349
rect 10749 23332 10754 23349
rect 10728 23328 10754 23332
rect 10820 23349 10846 23354
rect 10820 23332 10824 23349
rect 10824 23332 10841 23349
rect 10841 23332 10846 23349
rect 10820 23328 10846 23332
rect 6266 23315 6292 23320
rect 6266 23298 6270 23315
rect 6270 23298 6287 23315
rect 6287 23298 6292 23315
rect 6266 23294 6292 23298
rect 6634 23294 6660 23320
rect 9256 23294 9282 23320
rect 10406 23294 10432 23320
rect 6404 23281 6430 23286
rect 6404 23264 6408 23281
rect 6408 23264 6425 23281
rect 6425 23264 6430 23281
rect 6404 23260 6430 23264
rect 6726 23260 6752 23286
rect 9164 23260 9190 23286
rect 9348 23281 9374 23286
rect 9348 23264 9369 23281
rect 9369 23264 9374 23281
rect 9348 23260 9374 23264
rect 10636 23281 10662 23286
rect 10636 23264 10640 23281
rect 10640 23264 10657 23281
rect 10657 23264 10662 23281
rect 10636 23260 10662 23264
rect 10866 23260 10892 23286
rect 11648 23281 11674 23286
rect 11648 23264 11652 23281
rect 11652 23264 11669 23281
rect 11669 23264 11674 23281
rect 11648 23260 11674 23264
rect 6312 23247 6338 23252
rect 6312 23230 6316 23247
rect 6316 23230 6333 23247
rect 6333 23230 6338 23247
rect 6312 23226 6338 23230
rect 9026 23226 9052 23252
rect 12016 23315 12042 23320
rect 12016 23298 12020 23315
rect 12020 23298 12037 23315
rect 12037 23298 12042 23315
rect 12016 23294 12042 23298
rect 12108 23315 12134 23320
rect 12108 23298 12112 23315
rect 12112 23298 12129 23315
rect 12129 23298 12134 23315
rect 12108 23294 12134 23298
rect 14638 23349 14664 23354
rect 14638 23332 14642 23349
rect 14642 23332 14659 23349
rect 14659 23332 14664 23349
rect 14638 23328 14664 23332
rect 15236 23328 15262 23354
rect 17122 23349 17148 23354
rect 17122 23332 17126 23349
rect 17126 23332 17143 23349
rect 17143 23332 17148 23349
rect 17122 23328 17148 23332
rect 17950 23349 17976 23354
rect 17950 23332 17954 23349
rect 17954 23332 17971 23349
rect 17971 23332 17976 23349
rect 17950 23328 17976 23332
rect 12154 23281 12180 23286
rect 12154 23264 12158 23281
rect 12158 23264 12175 23281
rect 12175 23264 12180 23281
rect 12154 23260 12180 23264
rect 13120 23281 13146 23286
rect 13120 23264 13124 23281
rect 13124 23264 13141 23281
rect 13141 23264 13146 23281
rect 13120 23260 13146 23264
rect 13258 23281 13284 23286
rect 13258 23264 13262 23281
rect 13262 23264 13279 23281
rect 13279 23264 13284 23281
rect 14960 23294 14986 23320
rect 13258 23260 13284 23264
rect 12292 23226 12318 23252
rect 12844 23226 12870 23252
rect 14914 23260 14940 23286
rect 16294 23281 16320 23286
rect 16294 23264 16298 23281
rect 16298 23264 16315 23281
rect 16315 23264 16320 23281
rect 16294 23260 16320 23264
rect 16524 23281 16550 23286
rect 16524 23264 16528 23281
rect 16528 23264 16545 23281
rect 16545 23264 16550 23281
rect 17260 23294 17286 23320
rect 16524 23260 16550 23264
rect 15006 23226 15032 23252
rect 16570 23247 16596 23252
rect 16570 23230 16574 23247
rect 16574 23230 16591 23247
rect 16591 23230 16596 23247
rect 16570 23226 16596 23230
rect 17168 23260 17194 23286
rect 17904 23281 17930 23286
rect 17904 23264 17908 23281
rect 17908 23264 17925 23281
rect 17925 23264 17930 23281
rect 17904 23260 17930 23264
rect 18134 23281 18160 23286
rect 18134 23264 18138 23281
rect 18138 23264 18155 23281
rect 18155 23264 18160 23281
rect 18134 23260 18160 23264
rect 18502 23260 18528 23286
rect 19422 23260 19448 23286
rect 21216 23294 21242 23320
rect 21492 23315 21518 23320
rect 21492 23298 21509 23315
rect 21509 23298 21518 23315
rect 21492 23294 21518 23298
rect 21078 23260 21104 23286
rect 21354 23281 21380 23286
rect 21354 23264 21358 23281
rect 21358 23264 21375 23281
rect 21375 23264 21380 23281
rect 21354 23260 21380 23264
rect 16156 23192 16182 23218
rect 19376 23192 19402 23218
rect 6726 23158 6752 23184
rect 10406 23158 10432 23184
rect 12108 23158 12134 23184
rect 15236 23158 15262 23184
rect 21124 23179 21150 23184
rect 21124 23162 21128 23179
rect 21128 23162 21145 23179
rect 21145 23162 21150 23179
rect 21124 23158 21150 23162
rect 22044 23179 22070 23184
rect 22044 23162 22048 23179
rect 22048 23162 22065 23179
rect 22065 23162 22070 23179
rect 22044 23158 22070 23162
rect 6450 23056 6476 23082
rect 9532 23056 9558 23082
rect 6634 23022 6660 23048
rect 10866 23022 10892 23048
rect 4840 22988 4866 23014
rect 5162 22954 5188 22980
rect 5300 22954 5326 22980
rect 9256 22988 9282 23014
rect 12154 23056 12180 23082
rect 16524 23056 16550 23082
rect 17536 23077 17562 23082
rect 17536 23060 17540 23077
rect 17540 23060 17557 23077
rect 17557 23060 17562 23077
rect 17536 23056 17562 23060
rect 21262 23056 21288 23082
rect 21676 23077 21702 23082
rect 21676 23060 21680 23077
rect 21680 23060 21697 23077
rect 21697 23060 21702 23077
rect 21676 23056 21702 23060
rect 22688 23077 22714 23082
rect 22688 23060 22692 23077
rect 22692 23060 22709 23077
rect 22709 23060 22714 23077
rect 22688 23056 22714 23060
rect 14224 23022 14250 23048
rect 18410 23022 18436 23048
rect 18502 23022 18528 23048
rect 5254 22920 5280 22946
rect 5438 22920 5464 22946
rect 5530 22920 5556 22946
rect 5760 22920 5786 22946
rect 9394 22975 9420 22980
rect 9394 22958 9398 22975
rect 9398 22958 9415 22975
rect 9415 22958 9420 22975
rect 9394 22954 9420 22958
rect 11050 22954 11076 22980
rect 10268 22920 10294 22946
rect 14684 22988 14710 23014
rect 15098 23009 15124 23014
rect 15098 22992 15102 23009
rect 15102 22992 15119 23009
rect 15119 22992 15124 23009
rect 15098 22988 15124 22992
rect 17674 22988 17700 23014
rect 18548 22988 18574 23014
rect 19652 23009 19678 23014
rect 19652 22992 19656 23009
rect 19656 22992 19673 23009
rect 19673 22992 19678 23009
rect 19652 22988 19678 22992
rect 21078 23022 21104 23048
rect 21216 23009 21242 23014
rect 21216 22992 21220 23009
rect 21220 22992 21237 23009
rect 21237 22992 21242 23009
rect 21216 22988 21242 22992
rect 21308 22988 21334 23014
rect 11418 22954 11444 22980
rect 13120 22954 13146 22980
rect 13396 22954 13422 22980
rect 14500 22954 14526 22980
rect 14960 22975 14986 22980
rect 14960 22958 14964 22975
rect 14964 22958 14981 22975
rect 14981 22958 14986 22975
rect 14960 22954 14986 22958
rect 14408 22920 14434 22946
rect 16248 22975 16274 22980
rect 16248 22958 16252 22975
rect 16252 22958 16269 22975
rect 16269 22958 16274 22975
rect 16248 22954 16274 22958
rect 16524 22954 16550 22980
rect 16432 22920 16458 22946
rect 16708 22954 16734 22980
rect 17490 22975 17516 22980
rect 17490 22958 17494 22975
rect 17494 22958 17511 22975
rect 17511 22958 17516 22975
rect 17490 22954 17516 22958
rect 17582 22975 17608 22980
rect 17582 22958 17586 22975
rect 17586 22958 17603 22975
rect 17603 22958 17608 22975
rect 17582 22954 17608 22958
rect 17812 22975 17838 22980
rect 17812 22958 17816 22975
rect 17816 22958 17833 22975
rect 17833 22958 17838 22975
rect 17812 22954 17838 22958
rect 20158 22954 20184 22980
rect 20342 22975 20368 22980
rect 20342 22958 20346 22975
rect 20346 22958 20363 22975
rect 20363 22958 20368 22975
rect 20342 22954 20368 22958
rect 17398 22920 17424 22946
rect 17904 22920 17930 22946
rect 19790 22920 19816 22946
rect 21124 22954 21150 22980
rect 21584 22975 21610 22980
rect 21584 22958 21588 22975
rect 21588 22958 21605 22975
rect 21605 22958 21610 22975
rect 21584 22954 21610 22958
rect 21630 22975 21656 22980
rect 21630 22958 21634 22975
rect 21634 22958 21651 22975
rect 21651 22958 21656 22975
rect 21630 22954 21656 22958
rect 22044 22954 22070 22980
rect 22826 22954 22852 22980
rect 23194 22954 23220 22980
rect 24390 22954 24416 22980
rect 5944 22886 5970 22912
rect 9256 22886 9282 22912
rect 11556 22886 11582 22912
rect 16156 22886 16182 22912
rect 17950 22907 17976 22912
rect 17950 22890 17954 22907
rect 17954 22890 17971 22907
rect 17971 22890 17976 22907
rect 17950 22886 17976 22890
rect 20848 22886 20874 22912
rect 21216 22886 21242 22912
rect 24528 22920 24554 22946
rect 24850 22941 24876 22946
rect 24850 22924 24852 22941
rect 24852 22924 24876 22941
rect 24850 22920 24876 22924
rect 23378 22886 23404 22912
rect 25632 22886 25658 22912
rect 11648 22784 11674 22810
rect 14546 22784 14572 22810
rect 14684 22805 14710 22810
rect 14684 22788 14688 22805
rect 14688 22788 14705 22805
rect 14705 22788 14710 22805
rect 14684 22784 14710 22788
rect 14960 22784 14986 22810
rect 9716 22750 9742 22776
rect 3552 22737 3578 22742
rect 3552 22720 3573 22737
rect 3573 22720 3578 22737
rect 3552 22716 3578 22720
rect 3690 22716 3716 22742
rect 7324 22716 7350 22742
rect 7554 22716 7580 22742
rect 9348 22716 9374 22742
rect 11556 22716 11582 22742
rect 12982 22716 13008 22742
rect 13258 22716 13284 22742
rect 13718 22716 13744 22742
rect 3414 22703 3440 22708
rect 3414 22686 3418 22703
rect 3418 22686 3435 22703
rect 3435 22686 3440 22703
rect 3414 22682 3440 22686
rect 7278 22703 7304 22708
rect 7278 22686 7282 22703
rect 7282 22686 7299 22703
rect 7299 22686 7304 22703
rect 7278 22682 7304 22686
rect 9026 22682 9052 22708
rect 9670 22682 9696 22708
rect 14822 22716 14848 22742
rect 14960 22716 14986 22742
rect 17490 22750 17516 22776
rect 17812 22750 17838 22776
rect 19652 22784 19678 22810
rect 18548 22750 18574 22776
rect 21538 22750 21564 22776
rect 24850 22750 24876 22776
rect 28254 22750 28280 22776
rect 16248 22716 16274 22742
rect 17766 22737 17792 22742
rect 17766 22720 17783 22737
rect 17783 22720 17792 22737
rect 17766 22716 17792 22720
rect 17904 22716 17930 22742
rect 14914 22682 14940 22708
rect 15144 22682 15170 22708
rect 17628 22703 17654 22708
rect 17628 22686 17632 22703
rect 17632 22686 17649 22703
rect 17649 22686 17654 22703
rect 17628 22682 17654 22686
rect 18640 22682 18666 22708
rect 19606 22716 19632 22742
rect 21952 22716 21978 22742
rect 23286 22716 23312 22742
rect 28346 22737 28372 22742
rect 22090 22682 22116 22708
rect 13028 22648 13054 22674
rect 13626 22648 13652 22674
rect 19192 22648 19218 22674
rect 20158 22648 20184 22674
rect 4794 22614 4820 22640
rect 8658 22614 8684 22640
rect 17720 22614 17746 22640
rect 18502 22614 18528 22640
rect 18548 22614 18574 22640
rect 24160 22703 24186 22708
rect 24160 22686 24164 22703
rect 24164 22686 24181 22703
rect 24181 22686 24186 22703
rect 24160 22682 24186 22686
rect 28346 22720 28367 22737
rect 28367 22720 28372 22737
rect 28346 22716 28372 22720
rect 24252 22682 24278 22708
rect 28208 22703 28234 22708
rect 28208 22686 28212 22703
rect 28212 22686 28229 22703
rect 28229 22686 28234 22703
rect 28208 22682 28234 22686
rect 23332 22614 23358 22640
rect 24252 22635 24278 22640
rect 24252 22618 24256 22635
rect 24256 22618 24273 22635
rect 24273 22618 24278 22635
rect 24252 22614 24278 22618
rect 29726 22614 29752 22640
rect 6404 22512 6430 22538
rect 8290 22512 8316 22538
rect 17766 22512 17792 22538
rect 17904 22512 17930 22538
rect 23286 22533 23312 22538
rect 23286 22516 23290 22533
rect 23290 22516 23307 22533
rect 23307 22516 23312 22533
rect 23286 22512 23312 22516
rect 3138 22431 3164 22436
rect 3138 22414 3142 22431
rect 3142 22414 3159 22431
rect 3159 22414 3164 22431
rect 3138 22410 3164 22414
rect 3552 22410 3578 22436
rect 4840 22478 4866 22504
rect 4932 22478 4958 22504
rect 8658 22478 8684 22504
rect 4886 22444 4912 22470
rect 5024 22444 5050 22470
rect 7370 22444 7396 22470
rect 4794 22431 4820 22436
rect 4794 22414 4811 22431
rect 4811 22414 4820 22431
rect 4978 22431 5004 22436
rect 4794 22410 4820 22414
rect 3184 22376 3210 22402
rect 4978 22414 4989 22431
rect 4989 22414 5004 22431
rect 4978 22410 5004 22414
rect 5300 22431 5326 22436
rect 5300 22414 5304 22431
rect 5304 22414 5321 22431
rect 5321 22414 5326 22431
rect 5300 22410 5326 22414
rect 5576 22410 5602 22436
rect 5622 22410 5648 22436
rect 5944 22410 5970 22436
rect 7278 22410 7304 22436
rect 8336 22444 8362 22470
rect 16432 22478 16458 22504
rect 17628 22478 17654 22504
rect 23332 22478 23358 22504
rect 4656 22363 4682 22368
rect 4656 22346 4660 22363
rect 4660 22346 4677 22363
rect 4677 22346 4682 22363
rect 4656 22342 4682 22346
rect 4748 22342 4774 22368
rect 7462 22376 7488 22402
rect 7646 22397 7672 22402
rect 7646 22380 7648 22397
rect 7648 22380 7672 22397
rect 7646 22376 7672 22380
rect 8428 22376 8454 22402
rect 9072 22410 9098 22436
rect 13396 22431 13422 22436
rect 13396 22414 13400 22431
rect 13400 22414 13417 22431
rect 13417 22414 13422 22431
rect 13396 22410 13422 22414
rect 13718 22410 13744 22436
rect 14500 22410 14526 22436
rect 17674 22444 17700 22470
rect 18364 22444 18390 22470
rect 15052 22431 15078 22436
rect 15052 22414 15056 22431
rect 15056 22414 15073 22431
rect 15073 22414 15078 22431
rect 15052 22410 15078 22414
rect 16294 22431 16320 22436
rect 16294 22414 16298 22431
rect 16298 22414 16315 22431
rect 16315 22414 16320 22431
rect 16294 22410 16320 22414
rect 16616 22410 16642 22436
rect 17490 22410 17516 22436
rect 17950 22410 17976 22436
rect 21078 22410 21104 22436
rect 21354 22410 21380 22436
rect 21630 22410 21656 22436
rect 18502 22376 18528 22402
rect 21538 22397 21564 22402
rect 21538 22380 21540 22397
rect 21540 22380 21564 22397
rect 21538 22376 21564 22380
rect 23056 22431 23082 22436
rect 23056 22414 23060 22431
rect 23060 22414 23077 22431
rect 23077 22414 23082 22431
rect 23056 22410 23082 22414
rect 24252 22444 24278 22470
rect 24390 22465 24416 22470
rect 24390 22448 24394 22465
rect 24394 22448 24411 22465
rect 24411 22448 24416 22465
rect 24390 22444 24416 22448
rect 23378 22431 23404 22436
rect 23378 22414 23382 22431
rect 23382 22414 23399 22431
rect 23399 22414 23404 22431
rect 23378 22410 23404 22414
rect 24528 22431 24554 22436
rect 24528 22414 24549 22431
rect 24549 22414 24554 22431
rect 24528 22410 24554 22414
rect 24344 22376 24370 22402
rect 24436 22376 24462 22402
rect 26966 22410 26992 22436
rect 8980 22342 9006 22368
rect 13442 22363 13468 22368
rect 13442 22346 13446 22363
rect 13446 22346 13463 22363
rect 13463 22346 13468 22363
rect 13442 22342 13468 22346
rect 13856 22342 13882 22368
rect 13994 22342 14020 22368
rect 15236 22342 15262 22368
rect 15696 22342 15722 22368
rect 17582 22342 17608 22368
rect 17766 22342 17792 22368
rect 22734 22342 22760 22368
rect 23010 22363 23036 22368
rect 23010 22346 23014 22363
rect 23014 22346 23031 22363
rect 23031 22346 23036 22363
rect 23010 22342 23036 22346
rect 25402 22342 25428 22368
rect 4748 22240 4774 22266
rect 8428 22240 8454 22266
rect 9624 22240 9650 22266
rect 10360 22240 10386 22266
rect 14776 22240 14802 22266
rect 15144 22240 15170 22266
rect 18594 22240 18620 22266
rect 7002 22206 7028 22232
rect 9164 22206 9190 22232
rect 3552 22172 3578 22198
rect 3782 22172 3808 22198
rect 5208 22172 5234 22198
rect 7370 22193 7396 22198
rect 7370 22176 7391 22193
rect 7391 22176 7396 22193
rect 7370 22172 7396 22176
rect 9026 22172 9052 22198
rect 9808 22172 9834 22198
rect 14960 22193 14986 22198
rect 14960 22176 14964 22193
rect 14964 22176 14981 22193
rect 14981 22176 14986 22193
rect 14960 22172 14986 22176
rect 15052 22172 15078 22198
rect 16616 22206 16642 22232
rect 17168 22206 17194 22232
rect 17536 22206 17562 22232
rect 17904 22206 17930 22232
rect 3138 22138 3164 22164
rect 3414 22138 3440 22164
rect 7462 22070 7488 22096
rect 10314 22070 10340 22096
rect 17812 22172 17838 22198
rect 18548 22206 18574 22232
rect 21308 22227 21334 22232
rect 21308 22210 21310 22227
rect 21310 22210 21334 22227
rect 21308 22206 21334 22210
rect 23010 22206 23036 22232
rect 21078 22193 21104 22198
rect 21078 22176 21082 22193
rect 21082 22176 21099 22193
rect 21099 22176 21104 22193
rect 21078 22172 21104 22176
rect 21630 22172 21656 22198
rect 23332 22172 23358 22198
rect 24344 22227 24370 22232
rect 24344 22210 24348 22227
rect 24348 22210 24365 22227
rect 24365 22210 24370 22227
rect 24344 22206 24370 22210
rect 25632 22206 25658 22232
rect 25402 22193 25428 22198
rect 25402 22176 25406 22193
rect 25406 22176 25423 22193
rect 25423 22176 25428 22193
rect 25402 22172 25428 22176
rect 16432 22138 16458 22164
rect 17766 22159 17792 22164
rect 17766 22142 17770 22159
rect 17770 22142 17787 22159
rect 17787 22142 17792 22159
rect 17766 22138 17792 22142
rect 24206 22159 24232 22164
rect 24206 22142 24210 22159
rect 24210 22142 24227 22159
rect 24227 22142 24232 22159
rect 24206 22138 24232 22142
rect 24298 22138 24324 22164
rect 17398 22104 17424 22130
rect 18502 22125 18528 22130
rect 18502 22108 18506 22125
rect 18506 22108 18523 22125
rect 18523 22108 18528 22125
rect 18502 22104 18528 22108
rect 25586 22193 25612 22198
rect 25586 22176 25590 22193
rect 25590 22176 25607 22193
rect 25607 22176 25612 22193
rect 25586 22172 25612 22176
rect 26230 22206 26256 22232
rect 28530 22206 28556 22232
rect 26874 22172 26900 22198
rect 28208 22172 28234 22198
rect 28392 22193 28418 22198
rect 28392 22176 28413 22193
rect 28413 22176 28418 22193
rect 28392 22172 28418 22176
rect 26138 22138 26164 22164
rect 16708 22070 16734 22096
rect 22642 22070 22668 22096
rect 25678 22091 25704 22096
rect 25678 22074 25682 22091
rect 25682 22074 25699 22091
rect 25699 22074 25704 22091
rect 25678 22070 25704 22074
rect 27150 22070 27176 22096
rect 28024 22070 28050 22096
rect 29542 22070 29568 22096
rect 4932 21866 4958 21892
rect 5300 21968 5326 21994
rect 5346 21968 5372 21994
rect 5714 21968 5740 21994
rect 9716 21968 9742 21994
rect 5484 21866 5510 21892
rect 6450 21887 6476 21892
rect 6450 21870 6454 21887
rect 6454 21870 6471 21887
rect 6471 21870 6476 21887
rect 6450 21866 6476 21870
rect 6634 21900 6660 21926
rect 6726 21866 6752 21892
rect 10176 21887 10202 21892
rect 10176 21870 10180 21887
rect 10180 21870 10197 21887
rect 10197 21870 10202 21887
rect 10176 21866 10202 21870
rect 10268 21887 10294 21892
rect 10268 21870 10272 21887
rect 10272 21870 10289 21887
rect 10289 21870 10294 21887
rect 10268 21866 10294 21870
rect 10314 21887 10340 21892
rect 10314 21870 10318 21887
rect 10318 21870 10335 21887
rect 10335 21870 10340 21887
rect 10314 21866 10340 21870
rect 10360 21887 10386 21892
rect 10360 21870 10364 21887
rect 10364 21870 10381 21887
rect 10381 21870 10386 21887
rect 10360 21866 10386 21870
rect 11372 21866 11398 21892
rect 11464 21887 11490 21892
rect 11464 21870 11485 21887
rect 11485 21870 11490 21887
rect 11464 21866 11490 21870
rect 14500 21866 14526 21892
rect 5208 21832 5234 21858
rect 6634 21853 6660 21858
rect 6634 21836 6638 21853
rect 6638 21836 6655 21853
rect 6655 21836 6660 21853
rect 6634 21832 6660 21836
rect 11556 21853 11582 21858
rect 11556 21836 11558 21853
rect 11558 21836 11582 21853
rect 11556 21832 11582 21836
rect 14960 21887 14986 21892
rect 14960 21870 14964 21887
rect 14964 21870 14981 21887
rect 14981 21870 14986 21887
rect 14960 21866 14986 21870
rect 16616 21866 16642 21892
rect 17490 21968 17516 21994
rect 23056 21968 23082 21994
rect 17720 21900 17746 21926
rect 17904 21921 17930 21926
rect 17904 21904 17908 21921
rect 17908 21904 17925 21921
rect 17925 21904 17930 21921
rect 17904 21900 17930 21904
rect 19376 21900 19402 21926
rect 21078 21900 21104 21926
rect 17536 21887 17562 21892
rect 17536 21870 17540 21887
rect 17540 21870 17557 21887
rect 17557 21870 17562 21887
rect 17536 21866 17562 21870
rect 17812 21866 17838 21892
rect 19790 21866 19816 21892
rect 21124 21866 21150 21892
rect 21630 21866 21656 21892
rect 22504 21887 22530 21892
rect 22504 21870 22508 21887
rect 22508 21870 22525 21887
rect 22525 21870 22530 21887
rect 22504 21866 22530 21870
rect 22734 21900 22760 21926
rect 25586 21968 25612 21994
rect 26184 21968 26210 21994
rect 27380 21968 27406 21994
rect 25632 21934 25658 21960
rect 22642 21887 22668 21892
rect 22642 21870 22659 21887
rect 22659 21870 22668 21887
rect 22642 21866 22668 21870
rect 21446 21853 21472 21858
rect 21446 21836 21448 21853
rect 21448 21836 21472 21853
rect 21446 21832 21472 21836
rect 22320 21832 22346 21858
rect 23010 21866 23036 21892
rect 24390 21900 24416 21926
rect 23240 21887 23266 21892
rect 23240 21870 23244 21887
rect 23244 21870 23261 21887
rect 23261 21870 23266 21887
rect 23240 21866 23266 21870
rect 23332 21887 23358 21892
rect 6542 21819 6568 21824
rect 6542 21802 6546 21819
rect 6546 21802 6563 21819
rect 6563 21802 6568 21819
rect 6542 21798 6568 21802
rect 10590 21798 10616 21824
rect 12430 21798 12456 21824
rect 14086 21798 14112 21824
rect 14362 21798 14388 21824
rect 16340 21819 16366 21824
rect 16340 21802 16344 21819
rect 16344 21802 16361 21819
rect 16361 21802 16366 21819
rect 16340 21798 16366 21802
rect 16432 21798 16458 21824
rect 16524 21798 16550 21824
rect 20664 21798 20690 21824
rect 22504 21819 22530 21824
rect 22504 21802 22508 21819
rect 22508 21802 22525 21819
rect 22525 21802 22530 21819
rect 22504 21798 22530 21802
rect 23194 21832 23220 21858
rect 23332 21870 23336 21887
rect 23336 21870 23353 21887
rect 23353 21870 23358 21887
rect 23332 21866 23358 21870
rect 26230 21900 26256 21926
rect 25678 21866 25704 21892
rect 25862 21887 25888 21892
rect 25862 21870 25866 21887
rect 25866 21870 25883 21887
rect 25883 21870 25888 21887
rect 25862 21866 25888 21870
rect 26138 21866 26164 21892
rect 26874 21887 26900 21892
rect 26874 21870 26895 21887
rect 26895 21870 26900 21887
rect 26874 21866 26900 21870
rect 28024 21887 28050 21892
rect 28024 21870 28028 21887
rect 28028 21870 28045 21887
rect 28045 21870 28050 21887
rect 28024 21866 28050 21870
rect 28070 21887 28096 21892
rect 28070 21870 28085 21887
rect 28085 21870 28096 21887
rect 28070 21866 28096 21870
rect 28162 21887 28188 21892
rect 28162 21870 28186 21887
rect 28186 21870 28188 21887
rect 28162 21866 28188 21870
rect 28346 21887 28372 21892
rect 28346 21870 28357 21887
rect 28357 21870 28372 21887
rect 28346 21866 28372 21870
rect 24482 21832 24508 21858
rect 24666 21853 24692 21858
rect 24666 21836 24668 21853
rect 24668 21836 24692 21853
rect 24666 21832 24692 21836
rect 26966 21853 26992 21858
rect 26966 21836 26968 21853
rect 26968 21836 26992 21853
rect 26966 21832 26992 21836
rect 27196 21798 27222 21824
rect 6450 21696 6476 21722
rect 15512 21696 15538 21722
rect 3460 21662 3486 21688
rect 3644 21683 3670 21688
rect 3644 21666 3646 21683
rect 3646 21666 3670 21683
rect 3644 21662 3670 21666
rect 4656 21662 4682 21688
rect 7232 21662 7258 21688
rect 8520 21662 8546 21688
rect 9900 21683 9926 21688
rect 9900 21666 9902 21683
rect 9902 21666 9926 21683
rect 9900 21662 9926 21666
rect 11878 21683 11904 21688
rect 11878 21666 11880 21683
rect 11880 21666 11904 21683
rect 11878 21662 11904 21666
rect 12660 21662 12686 21688
rect 14546 21683 14572 21688
rect 14546 21666 14548 21683
rect 14548 21666 14572 21683
rect 14546 21662 14572 21666
rect 3552 21649 3578 21654
rect 3552 21632 3573 21649
rect 3573 21632 3578 21649
rect 3552 21628 3578 21632
rect 4840 21649 4866 21654
rect 4840 21632 4844 21649
rect 4844 21632 4861 21649
rect 4861 21632 4866 21649
rect 4840 21628 4866 21632
rect 4886 21649 4912 21654
rect 4886 21632 4890 21649
rect 4890 21632 4907 21649
rect 4907 21632 4912 21649
rect 4886 21628 4912 21632
rect 3414 21615 3440 21620
rect 3414 21598 3418 21615
rect 3418 21598 3435 21615
rect 3435 21598 3440 21615
rect 3414 21594 3440 21598
rect 6496 21649 6522 21654
rect 6496 21632 6500 21649
rect 6500 21632 6517 21649
rect 6517 21632 6522 21649
rect 6496 21628 6522 21632
rect 6542 21628 6568 21654
rect 7600 21628 7626 21654
rect 9670 21649 9696 21654
rect 9670 21632 9674 21649
rect 9674 21632 9691 21649
rect 9691 21632 9696 21649
rect 9670 21628 9696 21632
rect 9808 21649 9834 21654
rect 9808 21632 9829 21649
rect 9829 21632 9834 21649
rect 9808 21628 9834 21632
rect 11464 21628 11490 21654
rect 12706 21628 12732 21654
rect 13074 21649 13100 21654
rect 13074 21632 13078 21649
rect 13078 21632 13095 21649
rect 13095 21632 13100 21649
rect 13074 21628 13100 21632
rect 14224 21628 14250 21654
rect 15834 21649 15860 21654
rect 15834 21632 15838 21649
rect 15838 21632 15855 21649
rect 15855 21632 15860 21649
rect 15834 21628 15860 21632
rect 18226 21717 18252 21722
rect 18226 21700 18230 21717
rect 18230 21700 18247 21717
rect 18247 21700 18252 21717
rect 18226 21696 18252 21700
rect 21446 21696 21472 21722
rect 21676 21696 21702 21722
rect 22458 21696 22484 21722
rect 22550 21696 22576 21722
rect 25862 21696 25888 21722
rect 28162 21696 28188 21722
rect 16708 21662 16734 21688
rect 4702 21560 4728 21586
rect 4794 21526 4820 21552
rect 7278 21615 7304 21620
rect 7278 21598 7282 21615
rect 7282 21598 7299 21615
rect 7299 21598 7304 21615
rect 7278 21594 7304 21598
rect 11418 21594 11444 21620
rect 14178 21594 14204 21620
rect 16156 21649 16182 21654
rect 16156 21632 16160 21649
rect 16160 21632 16177 21649
rect 16177 21632 16182 21649
rect 16156 21628 16182 21632
rect 16248 21649 16274 21654
rect 16248 21632 16252 21649
rect 16252 21632 16269 21649
rect 16269 21632 16274 21649
rect 16248 21628 16274 21632
rect 17398 21628 17424 21654
rect 17720 21683 17746 21688
rect 17720 21666 17724 21683
rect 17724 21666 17741 21683
rect 17741 21666 17746 21683
rect 17720 21662 17746 21666
rect 16432 21594 16458 21620
rect 24666 21662 24692 21688
rect 26368 21683 26394 21688
rect 26368 21666 26370 21683
rect 26370 21666 26394 21683
rect 26368 21662 26394 21666
rect 28438 21683 28464 21688
rect 28438 21666 28440 21683
rect 28440 21666 28464 21683
rect 28438 21662 28464 21666
rect 26874 21628 26900 21654
rect 28208 21649 28234 21654
rect 28208 21632 28212 21649
rect 28212 21632 28229 21649
rect 28229 21632 28234 21649
rect 28208 21628 28234 21632
rect 28346 21649 28372 21654
rect 28346 21632 28367 21649
rect 28367 21632 28372 21649
rect 28346 21628 28372 21632
rect 29358 21628 29384 21654
rect 29542 21649 29568 21654
rect 29542 21632 29557 21649
rect 29557 21632 29568 21649
rect 29726 21662 29752 21688
rect 29542 21628 29568 21632
rect 29818 21649 29844 21654
rect 29818 21632 29829 21649
rect 29829 21632 29844 21649
rect 29818 21628 29844 21632
rect 17904 21594 17930 21620
rect 25540 21594 25566 21620
rect 26138 21615 26164 21620
rect 26138 21598 26142 21615
rect 26142 21598 26159 21615
rect 26159 21598 26164 21615
rect 26138 21594 26164 21598
rect 7646 21526 7672 21552
rect 8290 21526 8316 21552
rect 10774 21526 10800 21552
rect 12338 21526 12364 21552
rect 19468 21560 19494 21586
rect 29772 21560 29798 21586
rect 12614 21526 12640 21552
rect 29312 21526 29338 21552
rect 3690 21424 3716 21450
rect 4886 21390 4912 21416
rect 6634 21424 6660 21450
rect 7646 21424 7672 21450
rect 8520 21424 8546 21450
rect 8290 21390 8316 21416
rect 4932 21356 4958 21382
rect 9302 21424 9328 21450
rect 10176 21424 10202 21450
rect 5070 21322 5096 21348
rect 5346 21322 5372 21348
rect 5576 21322 5602 21348
rect 5714 21322 5740 21348
rect 4656 21309 4682 21314
rect 4656 21292 4660 21309
rect 4660 21292 4677 21309
rect 4677 21292 4682 21309
rect 4656 21288 4682 21292
rect 4748 21309 4774 21314
rect 4748 21292 4752 21309
rect 4752 21292 4769 21309
rect 4769 21292 4774 21309
rect 4748 21288 4774 21292
rect 4794 21309 4820 21314
rect 4794 21292 4798 21309
rect 4798 21292 4815 21309
rect 4815 21292 4820 21309
rect 4794 21288 4820 21292
rect 5530 21309 5556 21314
rect 5530 21292 5532 21309
rect 5532 21292 5556 21309
rect 5530 21288 5556 21292
rect 8244 21322 8270 21348
rect 8658 21343 8684 21348
rect 8658 21326 8662 21343
rect 8662 21326 8679 21343
rect 8679 21326 8684 21343
rect 8658 21322 8684 21326
rect 12982 21424 13008 21450
rect 16616 21445 16642 21450
rect 16616 21428 16620 21445
rect 16620 21428 16637 21445
rect 16637 21428 16642 21445
rect 16616 21424 16642 21428
rect 26184 21424 26210 21450
rect 29818 21424 29844 21450
rect 20388 21390 20414 21416
rect 24390 21390 24416 21416
rect 25540 21390 25566 21416
rect 9072 21322 9098 21348
rect 10590 21343 10616 21348
rect 10590 21326 10594 21343
rect 10594 21326 10611 21343
rect 10611 21326 10616 21343
rect 10590 21322 10616 21326
rect 10636 21343 10662 21348
rect 10636 21326 10640 21343
rect 10640 21326 10657 21343
rect 10657 21326 10662 21343
rect 10636 21322 10662 21326
rect 10774 21343 10800 21348
rect 10774 21326 10778 21343
rect 10778 21326 10795 21343
rect 10795 21326 10800 21343
rect 10774 21322 10800 21326
rect 10820 21343 10846 21348
rect 10820 21326 10824 21343
rect 10824 21326 10841 21343
rect 10841 21326 10846 21343
rect 10820 21322 10846 21326
rect 11050 21322 11076 21348
rect 11418 21343 11444 21348
rect 11418 21326 11422 21343
rect 11422 21326 11439 21343
rect 11439 21326 11444 21343
rect 11418 21322 11444 21326
rect 16248 21356 16274 21382
rect 19330 21377 19356 21382
rect 19330 21360 19334 21377
rect 19334 21360 19351 21377
rect 19351 21360 19356 21377
rect 19330 21356 19356 21360
rect 13074 21322 13100 21348
rect 14178 21343 14204 21348
rect 14178 21326 14182 21343
rect 14182 21326 14199 21343
rect 14199 21326 14204 21343
rect 14178 21322 14204 21326
rect 16708 21322 16734 21348
rect 17398 21322 17424 21348
rect 7278 21254 7304 21280
rect 7462 21254 7488 21280
rect 7968 21254 7994 21280
rect 8336 21254 8362 21280
rect 8888 21309 8914 21314
rect 8888 21292 8890 21309
rect 8890 21292 8914 21309
rect 8888 21288 8914 21292
rect 10866 21288 10892 21314
rect 10958 21288 10984 21314
rect 11464 21288 11490 21314
rect 11648 21309 11674 21314
rect 11648 21292 11650 21309
rect 11650 21292 11674 21309
rect 11648 21288 11674 21292
rect 13764 21288 13790 21314
rect 14224 21288 14250 21314
rect 14408 21309 14434 21314
rect 14408 21292 14410 21309
rect 14410 21292 14434 21309
rect 14408 21288 14434 21292
rect 19284 21288 19310 21314
rect 21216 21356 21242 21382
rect 21630 21356 21656 21382
rect 23700 21356 23726 21382
rect 24482 21356 24508 21382
rect 20342 21322 20368 21348
rect 24620 21322 24646 21348
rect 19560 21309 19586 21314
rect 19560 21292 19562 21309
rect 19562 21292 19586 21309
rect 19560 21288 19586 21292
rect 8612 21254 8638 21280
rect 8704 21254 8730 21280
rect 9670 21254 9696 21280
rect 10314 21254 10340 21280
rect 11050 21254 11076 21280
rect 12522 21254 12548 21280
rect 20112 21254 20138 21280
rect 24758 21288 24784 21314
rect 3552 21152 3578 21178
rect 6496 21173 6522 21178
rect 6496 21156 6500 21173
rect 6500 21156 6517 21173
rect 6517 21156 6522 21173
rect 6496 21152 6522 21156
rect 3184 21118 3210 21144
rect 3736 21139 3762 21144
rect 3414 21084 3440 21110
rect 3552 21084 3578 21110
rect 3736 21122 3738 21139
rect 3738 21122 3762 21139
rect 3736 21118 3762 21122
rect 4748 21118 4774 21144
rect 6588 21118 6614 21144
rect 6772 21118 6798 21144
rect 3920 21084 3946 21110
rect 4932 21105 4958 21110
rect 4932 21088 4936 21105
rect 4936 21088 4953 21105
rect 4953 21088 4958 21105
rect 4932 21084 4958 21088
rect 5208 21084 5234 21110
rect 5806 21084 5832 21110
rect 5116 21050 5142 21076
rect 4840 21016 4866 21042
rect 6542 21105 6568 21110
rect 6542 21088 6546 21105
rect 6546 21088 6563 21105
rect 6563 21088 6568 21105
rect 6542 21084 6568 21088
rect 6680 21105 6706 21110
rect 6680 21088 6684 21105
rect 6684 21088 6701 21105
rect 6701 21088 6706 21105
rect 6680 21084 6706 21088
rect 6818 21084 6844 21110
rect 8290 21152 8316 21178
rect 10636 21152 10662 21178
rect 12338 21152 12364 21178
rect 7232 21118 7258 21144
rect 7508 21139 7534 21144
rect 7508 21122 7510 21139
rect 7510 21122 7534 21139
rect 7508 21118 7534 21122
rect 9762 21139 9788 21144
rect 9762 21122 9764 21139
rect 9764 21122 9788 21139
rect 9762 21118 9788 21122
rect 12660 21152 12686 21178
rect 13074 21152 13100 21178
rect 16248 21152 16274 21178
rect 16386 21152 16412 21178
rect 20388 21152 20414 21178
rect 23884 21152 23910 21178
rect 7922 21084 7948 21110
rect 7968 21084 7994 21110
rect 8704 21084 8730 21110
rect 9808 21084 9834 21110
rect 10958 21084 10984 21110
rect 12384 21105 12410 21110
rect 12384 21088 12388 21105
rect 12388 21088 12405 21105
rect 12405 21088 12410 21105
rect 12384 21084 12410 21088
rect 12430 21105 12456 21110
rect 12430 21088 12445 21105
rect 12445 21088 12456 21105
rect 12430 21084 12456 21088
rect 12522 21105 12548 21110
rect 12522 21088 12546 21105
rect 12546 21088 12548 21105
rect 12522 21084 12548 21088
rect 12752 21084 12778 21110
rect 7278 21071 7304 21076
rect 7278 21054 7282 21071
rect 7282 21054 7299 21071
rect 7299 21054 7304 21071
rect 7278 21050 7304 21054
rect 8658 21050 8684 21076
rect 7922 20982 7948 21008
rect 9670 20982 9696 21008
rect 10222 20982 10248 21008
rect 11556 21050 11582 21076
rect 12614 21050 12640 21076
rect 12982 21118 13008 21144
rect 17260 21118 17286 21144
rect 18226 21118 18252 21144
rect 18548 21139 18574 21144
rect 18548 21122 18550 21139
rect 18550 21122 18574 21139
rect 18548 21118 18574 21122
rect 12936 21084 12962 21110
rect 16570 21084 16596 21110
rect 17214 21084 17240 21110
rect 20112 21105 20138 21110
rect 20112 21088 20116 21105
rect 20116 21088 20133 21105
rect 20133 21088 20138 21105
rect 20112 21084 20138 21088
rect 20342 21118 20368 21144
rect 20250 21105 20276 21110
rect 20250 21088 20267 21105
rect 20267 21088 20276 21105
rect 20480 21118 20506 21144
rect 20250 21084 20276 21088
rect 20940 21084 20966 21110
rect 23700 21084 23726 21110
rect 14270 21050 14296 21076
rect 14408 21050 14434 21076
rect 12660 21016 12686 21042
rect 16340 21016 16366 21042
rect 17168 21016 17194 21042
rect 19284 21050 19310 21076
rect 23378 21050 23404 21076
rect 19238 21016 19264 21042
rect 20388 21016 20414 21042
rect 20434 21016 20460 21042
rect 19008 20982 19034 21008
rect 19330 20982 19356 21008
rect 22642 20982 22668 21008
rect 23884 20982 23910 21008
rect 24574 20982 24600 21008
rect 25540 21084 25566 21110
rect 25724 21050 25750 21076
rect 26874 21084 26900 21110
rect 26368 20982 26394 21008
rect 27012 20982 27038 21008
rect 3414 20880 3440 20906
rect 4656 20880 4682 20906
rect 6680 20880 6706 20906
rect 7508 20880 7534 20906
rect 3552 20778 3578 20804
rect 5346 20778 5372 20804
rect 6956 20812 6982 20838
rect 7462 20812 7488 20838
rect 6726 20778 6752 20804
rect 6818 20778 6844 20804
rect 7554 20778 7580 20804
rect 8612 20880 8638 20906
rect 9578 20880 9604 20906
rect 11234 20880 11260 20906
rect 11280 20880 11306 20906
rect 11648 20880 11674 20906
rect 13074 20880 13100 20906
rect 12568 20846 12594 20872
rect 12798 20846 12824 20872
rect 10314 20812 10340 20838
rect 3184 20744 3210 20770
rect 3414 20744 3440 20770
rect 5760 20765 5786 20770
rect 5760 20748 5762 20765
rect 5762 20748 5786 20765
rect 5760 20744 5786 20748
rect 3920 20710 3946 20736
rect 5530 20710 5556 20736
rect 6358 20710 6384 20736
rect 7232 20710 7258 20736
rect 10958 20799 10984 20804
rect 10958 20782 10979 20799
rect 10979 20782 10984 20799
rect 10958 20778 10984 20782
rect 11832 20778 11858 20804
rect 12936 20812 12962 20838
rect 14178 20880 14204 20906
rect 17996 20880 18022 20906
rect 18548 20880 18574 20906
rect 20250 20880 20276 20906
rect 20434 20846 20460 20872
rect 19008 20833 19034 20838
rect 19008 20816 19012 20833
rect 19012 20816 19029 20833
rect 19029 20816 19034 20833
rect 19008 20812 19034 20816
rect 22504 20833 22530 20838
rect 22504 20816 22508 20833
rect 22508 20816 22525 20833
rect 22525 20816 22530 20833
rect 22504 20812 22530 20816
rect 24666 20833 24692 20838
rect 24666 20816 24670 20833
rect 24670 20816 24687 20833
rect 24687 20816 24692 20833
rect 24666 20812 24692 20816
rect 26874 20812 26900 20838
rect 28070 20880 28096 20906
rect 28208 20880 28234 20906
rect 13304 20778 13330 20804
rect 13028 20744 13054 20770
rect 19284 20778 19310 20804
rect 21078 20778 21104 20804
rect 22642 20799 22668 20804
rect 22642 20782 22646 20799
rect 22646 20782 22663 20799
rect 22663 20782 22668 20799
rect 22642 20778 22668 20782
rect 24758 20799 24784 20804
rect 24758 20782 24765 20799
rect 24765 20782 24782 20799
rect 24782 20782 24784 20799
rect 24758 20778 24784 20782
rect 27058 20778 27084 20804
rect 28116 20799 28142 20804
rect 28116 20782 28137 20799
rect 28137 20782 28142 20799
rect 28116 20778 28142 20782
rect 28254 20778 28280 20804
rect 11280 20710 11306 20736
rect 12614 20710 12640 20736
rect 13074 20710 13100 20736
rect 13764 20744 13790 20770
rect 19238 20765 19264 20770
rect 19238 20748 19240 20765
rect 19240 20748 19264 20765
rect 19238 20744 19264 20748
rect 21446 20765 21472 20770
rect 21446 20748 21448 20765
rect 21448 20748 21472 20765
rect 21446 20744 21472 20748
rect 22688 20765 22714 20770
rect 22688 20748 22692 20765
rect 22692 20748 22709 20765
rect 22709 20748 22714 20765
rect 22688 20744 22714 20748
rect 22872 20765 22898 20770
rect 22872 20748 22876 20765
rect 22876 20748 22893 20765
rect 22893 20748 22898 20765
rect 22872 20744 22898 20748
rect 24574 20765 24600 20770
rect 24574 20748 24578 20765
rect 24578 20748 24595 20765
rect 24595 20748 24600 20765
rect 24574 20744 24600 20748
rect 24620 20744 24646 20770
rect 14868 20710 14894 20736
rect 21216 20710 21242 20736
rect 22550 20710 22576 20736
rect 22596 20731 22622 20736
rect 22596 20714 22600 20731
rect 22600 20714 22617 20731
rect 22617 20714 22622 20731
rect 22596 20710 22622 20714
rect 24712 20765 24738 20770
rect 24712 20748 24716 20765
rect 24716 20748 24733 20765
rect 24733 20748 24738 20765
rect 24712 20744 24738 20748
rect 27196 20710 27222 20736
rect 29588 20710 29614 20736
rect 4932 20608 4958 20634
rect 5530 20608 5556 20634
rect 5714 20608 5740 20634
rect 3828 20574 3854 20600
rect 7922 20629 7948 20634
rect 7922 20612 7926 20629
rect 7926 20612 7943 20629
rect 7943 20612 7948 20629
rect 7922 20608 7948 20612
rect 15512 20629 15538 20634
rect 15512 20612 15516 20629
rect 15516 20612 15533 20629
rect 15533 20612 15538 20629
rect 15512 20608 15538 20612
rect 24712 20608 24738 20634
rect 29588 20608 29614 20634
rect 3552 20540 3578 20566
rect 3920 20561 3946 20566
rect 3920 20544 3941 20561
rect 3941 20544 3946 20561
rect 6358 20574 6384 20600
rect 7600 20574 7626 20600
rect 3920 20540 3946 20544
rect 4472 20540 4498 20566
rect 6496 20561 6522 20566
rect 6496 20544 6517 20561
rect 6517 20544 6522 20561
rect 6496 20540 6522 20544
rect 7002 20540 7028 20566
rect 7692 20540 7718 20566
rect 7784 20561 7810 20566
rect 7784 20544 7788 20561
rect 7788 20544 7805 20561
rect 7805 20544 7810 20561
rect 7784 20540 7810 20544
rect 7830 20561 7856 20566
rect 7830 20544 7834 20561
rect 7834 20544 7851 20561
rect 7851 20544 7856 20561
rect 7830 20540 7856 20544
rect 8290 20540 8316 20566
rect 11372 20540 11398 20566
rect 11464 20540 11490 20566
rect 14224 20574 14250 20600
rect 21124 20574 21150 20600
rect 6174 20506 6200 20532
rect 10268 20506 10294 20532
rect 11050 20506 11076 20532
rect 11418 20506 11444 20532
rect 7646 20472 7672 20498
rect 7692 20472 7718 20498
rect 8980 20472 9006 20498
rect 10176 20472 10202 20498
rect 14776 20561 14802 20566
rect 14776 20544 14780 20561
rect 14780 20544 14797 20561
rect 14797 20544 14802 20561
rect 14776 20540 14802 20544
rect 14868 20561 14894 20566
rect 14868 20544 14872 20561
rect 14872 20544 14889 20561
rect 14889 20544 14894 20561
rect 14868 20540 14894 20544
rect 15282 20561 15308 20566
rect 15282 20544 15286 20561
rect 15286 20544 15303 20561
rect 15303 20544 15308 20561
rect 15282 20540 15308 20544
rect 12798 20506 12824 20532
rect 13028 20506 13054 20532
rect 15374 20561 15400 20566
rect 15374 20544 15378 20561
rect 15378 20544 15395 20561
rect 15395 20544 15400 20561
rect 15374 20540 15400 20544
rect 21216 20540 21242 20566
rect 21354 20540 21380 20566
rect 22550 20574 22576 20600
rect 21078 20527 21104 20532
rect 21078 20510 21082 20527
rect 21082 20510 21099 20527
rect 21099 20510 21104 20527
rect 21078 20506 21104 20510
rect 15006 20472 15032 20498
rect 12384 20438 12410 20464
rect 13028 20438 13054 20464
rect 13442 20438 13468 20464
rect 15926 20438 15952 20464
rect 17030 20438 17056 20464
rect 22642 20540 22668 20566
rect 22918 20540 22944 20566
rect 23562 20540 23588 20566
rect 23654 20561 23680 20566
rect 23654 20544 23675 20561
rect 23675 20544 23680 20561
rect 25586 20574 25612 20600
rect 28116 20574 28142 20600
rect 23654 20540 23680 20544
rect 23930 20540 23956 20566
rect 25678 20561 25704 20566
rect 25678 20544 25699 20561
rect 25699 20544 25704 20561
rect 25678 20540 25704 20544
rect 26828 20561 26854 20566
rect 26828 20544 26832 20561
rect 26832 20544 26849 20561
rect 26849 20544 26854 20561
rect 26828 20540 26854 20544
rect 23056 20506 23082 20532
rect 23378 20506 23404 20532
rect 25540 20527 25566 20532
rect 25540 20510 25544 20527
rect 25544 20510 25561 20527
rect 25561 20510 25566 20527
rect 25540 20506 25566 20510
rect 22688 20472 22714 20498
rect 23240 20438 23266 20464
rect 26230 20438 26256 20464
rect 26782 20438 26808 20464
rect 28530 20540 28556 20566
rect 29358 20540 29384 20566
rect 29542 20561 29568 20566
rect 29542 20544 29559 20561
rect 29559 20544 29568 20561
rect 29542 20540 29568 20544
rect 28070 20506 28096 20532
rect 29266 20506 29292 20532
rect 29818 20540 29844 20566
rect 29772 20506 29798 20532
rect 5530 20336 5556 20362
rect 6542 20336 6568 20362
rect 9026 20336 9052 20362
rect 11878 20336 11904 20362
rect 12016 20336 12042 20362
rect 12752 20336 12778 20362
rect 14224 20357 14250 20362
rect 14224 20340 14228 20357
rect 14228 20340 14245 20357
rect 14245 20340 14250 20357
rect 14224 20336 14250 20340
rect 15374 20336 15400 20362
rect 19376 20336 19402 20362
rect 19790 20336 19816 20362
rect 21446 20336 21472 20362
rect 25586 20336 25612 20362
rect 26828 20336 26854 20362
rect 28254 20336 28280 20362
rect 28438 20336 28464 20362
rect 29542 20336 29568 20362
rect 3552 20234 3578 20260
rect 5346 20255 5372 20260
rect 5346 20238 5350 20255
rect 5350 20238 5367 20255
rect 5367 20238 5372 20255
rect 5346 20234 5372 20238
rect 11418 20289 11444 20294
rect 11418 20272 11422 20289
rect 11422 20272 11439 20289
rect 11439 20272 11444 20289
rect 11418 20268 11444 20272
rect 12752 20268 12778 20294
rect 12936 20289 12962 20294
rect 12936 20272 12940 20289
rect 12940 20272 12957 20289
rect 12957 20272 12962 20289
rect 12936 20268 12962 20272
rect 5760 20234 5786 20260
rect 6082 20234 6108 20260
rect 10406 20234 10432 20260
rect 11142 20234 11168 20260
rect 12798 20234 12824 20260
rect 13074 20255 13100 20260
rect 13074 20238 13095 20255
rect 13095 20238 13100 20255
rect 13074 20234 13100 20238
rect 13626 20234 13652 20260
rect 14316 20255 14342 20260
rect 14316 20238 14322 20255
rect 14322 20238 14342 20255
rect 14316 20234 14342 20238
rect 11372 20200 11398 20226
rect 13166 20221 13192 20226
rect 13166 20204 13168 20221
rect 13168 20204 13192 20221
rect 13166 20200 13192 20204
rect 6404 20166 6430 20192
rect 7048 20166 7074 20192
rect 9026 20166 9052 20192
rect 12430 20166 12456 20192
rect 14224 20166 14250 20192
rect 14423 20255 14449 20260
rect 14423 20238 14427 20255
rect 14427 20238 14444 20255
rect 14444 20238 14449 20255
rect 14423 20234 14449 20238
rect 14362 20166 14388 20192
rect 14423 20166 14449 20192
rect 14730 20234 14756 20260
rect 15098 20234 15124 20260
rect 27012 20302 27038 20328
rect 15880 20268 15906 20294
rect 16892 20268 16918 20294
rect 17168 20268 17194 20294
rect 15190 20234 15216 20260
rect 15420 20234 15446 20260
rect 17214 20234 17240 20260
rect 17306 20255 17332 20260
rect 17306 20238 17321 20255
rect 17321 20238 17332 20255
rect 17306 20234 17332 20238
rect 17398 20255 17424 20260
rect 19330 20268 19356 20294
rect 17398 20238 17422 20255
rect 17422 20238 17424 20255
rect 17398 20234 17424 20238
rect 15282 20200 15308 20226
rect 15834 20200 15860 20226
rect 15926 20166 15952 20192
rect 15972 20166 15998 20192
rect 17076 20166 17102 20192
rect 19560 20234 19586 20260
rect 19376 20200 19402 20226
rect 20894 20234 20920 20260
rect 22642 20234 22668 20260
rect 26322 20234 26348 20260
rect 26782 20255 26808 20260
rect 26782 20238 26797 20255
rect 26797 20238 26808 20255
rect 26782 20234 26808 20238
rect 27058 20255 27084 20260
rect 27058 20238 27069 20255
rect 27069 20238 27084 20255
rect 27058 20234 27084 20238
rect 28024 20234 28050 20260
rect 28116 20255 28142 20260
rect 28116 20238 28137 20255
rect 28137 20238 28142 20255
rect 28116 20234 28142 20238
rect 28300 20234 28326 20260
rect 27334 20200 27360 20226
rect 27794 20200 27820 20226
rect 28254 20200 28280 20226
rect 20802 20166 20828 20192
rect 23286 20166 23312 20192
rect 24114 20166 24140 20192
rect 26920 20166 26946 20192
rect 10268 20064 10294 20090
rect 12016 20064 12042 20090
rect 12430 20064 12456 20090
rect 14362 20064 14388 20090
rect 18364 20064 18390 20090
rect 19238 20064 19264 20090
rect 6404 20051 6430 20056
rect 6404 20034 6406 20051
rect 6406 20034 6430 20051
rect 6404 20030 6430 20034
rect 9026 20051 9052 20056
rect 9026 20034 9028 20051
rect 9028 20034 9052 20051
rect 9026 20030 9052 20034
rect 10176 20051 10202 20056
rect 10176 20034 10180 20051
rect 10180 20034 10197 20051
rect 10197 20034 10202 20051
rect 10176 20030 10202 20034
rect 6496 19996 6522 20022
rect 7784 19996 7810 20022
rect 8658 19996 8684 20022
rect 9072 19996 9098 20022
rect 9348 19996 9374 20022
rect 10084 20017 10110 20022
rect 10084 20000 10088 20017
rect 10088 20000 10105 20017
rect 10105 20000 10110 20017
rect 10084 19996 10110 20000
rect 5668 19962 5694 19988
rect 6174 19983 6200 19988
rect 6174 19966 6178 19983
rect 6178 19966 6195 19983
rect 6195 19966 6200 19983
rect 6174 19962 6200 19966
rect 10268 20017 10294 20022
rect 10268 20000 10275 20017
rect 10275 20000 10292 20017
rect 10292 20000 10294 20017
rect 10268 19996 10294 20000
rect 11786 19996 11812 20022
rect 11878 20017 11904 20022
rect 11878 20000 11882 20017
rect 11882 20000 11899 20017
rect 11899 20000 11904 20017
rect 11878 19996 11904 20000
rect 11924 20017 11950 20022
rect 11924 20000 11928 20017
rect 11928 20000 11945 20017
rect 11945 20000 11950 20017
rect 11924 19996 11950 20000
rect 12338 19996 12364 20022
rect 12384 20017 12410 20022
rect 12384 20000 12388 20017
rect 12388 20000 12405 20017
rect 12405 20000 12410 20017
rect 12384 19996 12410 20000
rect 12614 20030 12640 20056
rect 13028 20051 13054 20056
rect 13028 20034 13030 20051
rect 13030 20034 13054 20051
rect 13028 20030 13054 20034
rect 15604 20030 15630 20056
rect 13120 19996 13146 20022
rect 15006 19996 15032 20022
rect 15144 19996 15170 20022
rect 15972 19996 15998 20022
rect 16110 19996 16136 20022
rect 17306 19996 17332 20022
rect 17858 20017 17884 20022
rect 17858 20000 17879 20017
rect 17879 20000 17884 20017
rect 17858 19996 17884 20000
rect 18364 19996 18390 20022
rect 20802 20051 20828 20056
rect 20802 20034 20806 20051
rect 20806 20034 20823 20051
rect 20823 20034 20828 20051
rect 20802 20030 20828 20034
rect 23286 20030 23312 20056
rect 24114 20030 24140 20056
rect 12614 19962 12640 19988
rect 12752 19962 12778 19988
rect 9348 19894 9374 19920
rect 10314 19894 10340 19920
rect 12706 19928 12732 19954
rect 12062 19894 12088 19920
rect 17720 19983 17746 19988
rect 17720 19966 17724 19983
rect 17724 19966 17741 19983
rect 17741 19966 17746 19983
rect 17720 19962 17746 19966
rect 20342 19996 20368 20022
rect 20572 19996 20598 20022
rect 20664 20017 20690 20022
rect 20664 20000 20668 20017
rect 20668 20000 20685 20017
rect 20685 20000 20690 20017
rect 20664 19996 20690 20000
rect 20756 20017 20782 20022
rect 20756 20000 20760 20017
rect 20760 20000 20777 20017
rect 20777 20000 20782 20017
rect 20756 19996 20782 20000
rect 20940 19996 20966 20022
rect 22688 19996 22714 20022
rect 23056 19996 23082 20022
rect 23148 20017 23174 20022
rect 23148 20000 23169 20017
rect 23169 20000 23174 20017
rect 23148 19996 23174 20000
rect 23562 19996 23588 20022
rect 24436 20017 24462 20022
rect 24436 20000 24440 20017
rect 24440 20000 24457 20017
rect 24457 20000 24462 20017
rect 24436 19996 24462 20000
rect 24482 20017 24508 20022
rect 24482 20000 24489 20017
rect 24489 20000 24506 20017
rect 24506 20000 24508 20017
rect 24482 19996 24508 20000
rect 25540 19996 25566 20022
rect 25724 20017 25750 20022
rect 25724 20000 25745 20017
rect 25745 20000 25750 20017
rect 25724 19996 25750 20000
rect 26920 19996 26946 20022
rect 20894 19928 20920 19954
rect 22964 19928 22990 19954
rect 15880 19894 15906 19920
rect 15972 19894 15998 19920
rect 18870 19894 18896 19920
rect 20664 19894 20690 19920
rect 23102 19894 23128 19920
rect 24252 19894 24278 19920
rect 24298 19915 24324 19920
rect 24298 19898 24302 19915
rect 24302 19898 24319 19915
rect 24319 19898 24324 19915
rect 24298 19894 24324 19898
rect 24482 19894 24508 19920
rect 29266 19894 29292 19920
rect 5346 19724 5372 19750
rect 5668 19792 5694 19818
rect 10084 19792 10110 19818
rect 8658 19745 8684 19750
rect 8658 19728 8662 19745
rect 8662 19728 8679 19745
rect 8679 19728 8684 19745
rect 8658 19724 8684 19728
rect 9578 19724 9604 19750
rect 10728 19724 10754 19750
rect 11050 19792 11076 19818
rect 11878 19792 11904 19818
rect 12062 19792 12088 19818
rect 12522 19758 12548 19784
rect 12614 19758 12640 19784
rect 14362 19792 14388 19818
rect 17398 19792 17424 19818
rect 14730 19758 14756 19784
rect 19330 19724 19356 19750
rect 5530 19711 5556 19716
rect 5530 19694 5551 19711
rect 5551 19694 5556 19711
rect 5530 19690 5556 19694
rect 9072 19690 9098 19716
rect 10314 19711 10340 19716
rect 10314 19694 10318 19711
rect 10318 19694 10335 19711
rect 10335 19694 10340 19711
rect 10314 19690 10340 19694
rect 10360 19711 10386 19716
rect 10360 19694 10364 19711
rect 10364 19694 10381 19711
rect 10381 19694 10386 19711
rect 10360 19690 10386 19694
rect 11372 19690 11398 19716
rect 12752 19690 12778 19716
rect 13028 19690 13054 19716
rect 13304 19690 13330 19716
rect 15972 19711 15998 19716
rect 15972 19694 15976 19711
rect 15976 19694 15993 19711
rect 15993 19694 15998 19711
rect 15972 19690 15998 19694
rect 16110 19711 16136 19716
rect 16110 19694 16131 19711
rect 16131 19694 16136 19711
rect 21446 19792 21472 19818
rect 24252 19792 24278 19818
rect 27334 19792 27360 19818
rect 22688 19758 22714 19784
rect 24482 19758 24508 19784
rect 16110 19690 16136 19694
rect 5622 19677 5648 19682
rect 5622 19660 5624 19677
rect 5624 19660 5648 19677
rect 5622 19656 5648 19660
rect 8704 19656 8730 19682
rect 11188 19677 11214 19682
rect 11188 19660 11190 19677
rect 11190 19660 11214 19677
rect 11188 19656 11214 19660
rect 16248 19656 16274 19682
rect 19376 19656 19402 19682
rect 21078 19690 21104 19716
rect 21262 19690 21288 19716
rect 21584 19690 21610 19716
rect 23286 19690 23312 19716
rect 21354 19656 21380 19682
rect 6404 19622 6430 19648
rect 12982 19622 13008 19648
rect 20434 19622 20460 19648
rect 22734 19622 22760 19648
rect 22964 19622 22990 19648
rect 27794 19622 27820 19648
rect 11188 19520 11214 19546
rect 12614 19520 12640 19546
rect 13166 19520 13192 19546
rect 20572 19541 20598 19546
rect 20572 19524 20576 19541
rect 20576 19524 20593 19541
rect 20593 19524 20598 19541
rect 20572 19520 20598 19524
rect 22596 19541 22622 19546
rect 22596 19524 22600 19541
rect 22600 19524 22617 19541
rect 22617 19524 22622 19541
rect 22596 19520 22622 19524
rect 22780 19520 22806 19546
rect 3782 19507 3808 19512
rect 3782 19490 3784 19507
rect 3784 19490 3808 19507
rect 3782 19486 3808 19490
rect 4978 19486 5004 19512
rect 3552 19473 3578 19478
rect 3552 19456 3556 19473
rect 3556 19456 3573 19473
rect 3573 19456 3578 19473
rect 3552 19452 3578 19456
rect 3598 19452 3624 19478
rect 4840 19473 4866 19478
rect 4840 19456 4844 19473
rect 4844 19456 4861 19473
rect 4861 19456 4866 19473
rect 4840 19452 4866 19456
rect 4932 19473 4958 19478
rect 4932 19456 4938 19473
rect 4938 19456 4958 19473
rect 4932 19452 4958 19456
rect 7554 19486 7580 19512
rect 5162 19473 5188 19478
rect 5162 19456 5173 19473
rect 5173 19456 5188 19473
rect 4932 19384 4958 19410
rect 5024 19418 5050 19444
rect 4840 19371 4866 19376
rect 4840 19354 4844 19371
rect 4844 19354 4861 19371
rect 4861 19354 4866 19371
rect 4840 19350 4866 19354
rect 5162 19452 5188 19456
rect 7278 19473 7304 19478
rect 7278 19456 7282 19473
rect 7282 19456 7299 19473
rect 7299 19456 7304 19473
rect 7278 19452 7304 19456
rect 7416 19473 7442 19478
rect 7416 19456 7437 19473
rect 7437 19456 7442 19473
rect 7416 19452 7442 19456
rect 8382 19452 8408 19478
rect 8842 19473 8868 19478
rect 20066 19486 20092 19512
rect 20434 19507 20460 19512
rect 20434 19490 20438 19507
rect 20438 19490 20455 19507
rect 20455 19490 20460 19507
rect 20434 19486 20460 19490
rect 21308 19507 21334 19512
rect 21308 19490 21310 19507
rect 21310 19490 21334 19507
rect 21308 19486 21334 19490
rect 24436 19520 24462 19546
rect 22964 19486 22990 19512
rect 8842 19456 8857 19473
rect 8857 19456 8868 19473
rect 8842 19452 8868 19456
rect 9118 19473 9144 19478
rect 9118 19456 9129 19473
rect 9129 19456 9144 19473
rect 8244 19384 8270 19410
rect 9118 19452 9144 19456
rect 9210 19452 9236 19478
rect 12522 19452 12548 19478
rect 20296 19473 20322 19478
rect 20296 19456 20300 19473
rect 20300 19456 20317 19473
rect 20317 19456 20322 19473
rect 20296 19452 20322 19456
rect 9302 19418 9328 19444
rect 9624 19418 9650 19444
rect 8980 19384 9006 19410
rect 9302 19350 9328 19376
rect 12384 19350 12410 19376
rect 21032 19452 21058 19478
rect 21354 19452 21380 19478
rect 22596 19473 22622 19478
rect 22596 19456 22600 19473
rect 22600 19456 22617 19473
rect 22617 19456 22622 19473
rect 22596 19452 22622 19456
rect 21078 19439 21104 19444
rect 21078 19422 21082 19439
rect 21082 19422 21099 19439
rect 21099 19422 21104 19439
rect 21078 19418 21104 19422
rect 22734 19473 22760 19478
rect 22734 19456 22751 19473
rect 22751 19456 22760 19473
rect 22734 19452 22760 19456
rect 22918 19473 22944 19478
rect 22918 19456 22929 19473
rect 22929 19456 22944 19473
rect 22918 19452 22944 19456
rect 23194 19452 23220 19478
rect 22964 19418 22990 19444
rect 23056 19418 23082 19444
rect 22642 19350 22668 19376
rect 22826 19350 22852 19376
rect 23102 19350 23128 19376
rect 4886 19248 4912 19274
rect 5668 19248 5694 19274
rect 5806 19248 5832 19274
rect 3138 19167 3164 19172
rect 3138 19150 3142 19167
rect 3142 19150 3159 19167
rect 3159 19150 3164 19167
rect 3138 19146 3164 19150
rect 3552 19146 3578 19172
rect 5576 19146 5602 19172
rect 8244 19248 8270 19274
rect 8842 19248 8868 19274
rect 17720 19248 17746 19274
rect 7278 19180 7304 19206
rect 19238 19248 19264 19274
rect 19330 19248 19356 19274
rect 20296 19248 20322 19274
rect 22780 19248 22806 19274
rect 25540 19248 25566 19274
rect 25632 19248 25658 19274
rect 26690 19214 26716 19240
rect 20710 19180 20736 19206
rect 3368 19133 3394 19138
rect 3368 19116 3370 19133
rect 3370 19116 3394 19133
rect 3368 19112 3394 19116
rect 8290 19146 8316 19172
rect 8474 19146 8500 19172
rect 18640 19146 18666 19172
rect 21262 19146 21288 19172
rect 21354 19146 21380 19172
rect 27380 19201 27406 19206
rect 27380 19184 27384 19201
rect 27384 19184 27401 19201
rect 27401 19184 27406 19201
rect 27380 19180 27406 19184
rect 6818 19133 6844 19138
rect 6818 19116 6822 19133
rect 6822 19116 6839 19133
rect 6839 19116 6844 19133
rect 6818 19112 6844 19116
rect 6910 19133 6936 19138
rect 6910 19116 6914 19133
rect 6914 19116 6931 19133
rect 6931 19116 6936 19133
rect 6910 19112 6936 19116
rect 7416 19112 7442 19138
rect 5576 19078 5602 19104
rect 6542 19078 6568 19104
rect 12108 19078 12134 19104
rect 12982 19078 13008 19104
rect 17950 19078 17976 19104
rect 21032 19112 21058 19138
rect 24160 19078 24186 19104
rect 24436 19112 24462 19138
rect 29542 19146 29568 19172
rect 28622 19112 28648 19138
rect 25494 19078 25520 19104
rect 27242 19099 27268 19104
rect 27242 19082 27246 19099
rect 27246 19082 27263 19099
rect 27263 19082 27268 19099
rect 27242 19078 27268 19082
rect 27288 19099 27314 19104
rect 27288 19082 27292 19099
rect 27292 19082 27309 19099
rect 27309 19082 27314 19099
rect 27288 19078 27314 19082
rect 4840 18976 4866 19002
rect 6818 18976 6844 19002
rect 8980 18976 9006 19002
rect 14960 18976 14986 19002
rect 3690 18942 3716 18968
rect 6496 18963 6522 18968
rect 6496 18946 6500 18963
rect 6500 18946 6517 18963
rect 6517 18946 6522 18963
rect 6496 18942 6522 18946
rect 6542 18963 6568 18968
rect 6542 18946 6546 18963
rect 6546 18946 6563 18963
rect 6563 18946 6568 18963
rect 6542 18942 6568 18946
rect 7508 18963 7534 18968
rect 7508 18946 7510 18963
rect 7510 18946 7534 18963
rect 7508 18942 7534 18946
rect 3138 18908 3164 18934
rect 3552 18929 3578 18934
rect 3552 18912 3573 18929
rect 3573 18912 3578 18929
rect 3552 18908 3578 18912
rect 4702 18874 4728 18900
rect 4840 18929 4866 18934
rect 4840 18912 4844 18929
rect 4844 18912 4861 18929
rect 4861 18912 4866 18929
rect 4840 18908 4866 18912
rect 6404 18929 6430 18934
rect 6404 18912 6408 18929
rect 6408 18912 6425 18929
rect 6425 18912 6430 18929
rect 6404 18908 6430 18912
rect 6634 18908 6660 18934
rect 7278 18929 7304 18934
rect 7278 18912 7282 18929
rect 7282 18912 7299 18929
rect 7299 18912 7304 18929
rect 7278 18908 7304 18912
rect 7416 18929 7442 18934
rect 6956 18874 6982 18900
rect 7416 18912 7437 18929
rect 7437 18912 7442 18929
rect 7416 18908 7442 18912
rect 11464 18908 11490 18934
rect 12108 18908 12134 18934
rect 14316 18942 14342 18968
rect 24298 18976 24324 19002
rect 24666 18976 24692 19002
rect 12430 18908 12456 18934
rect 12568 18908 12594 18934
rect 14592 18908 14618 18934
rect 15052 18908 15078 18934
rect 15696 18929 15722 18934
rect 15696 18912 15700 18929
rect 15700 18912 15717 18929
rect 15717 18912 15722 18929
rect 15696 18908 15722 18912
rect 15742 18929 15768 18934
rect 15742 18912 15746 18929
rect 15746 18912 15763 18929
rect 15763 18912 15768 18929
rect 15742 18908 15768 18912
rect 11832 18895 11858 18900
rect 11832 18878 11836 18895
rect 11836 18878 11853 18895
rect 11853 18878 11858 18895
rect 11832 18874 11858 18878
rect 14086 18874 14112 18900
rect 15282 18874 15308 18900
rect 15650 18874 15676 18900
rect 17720 18908 17746 18934
rect 17950 18908 17976 18934
rect 21354 18942 21380 18968
rect 22964 18942 22990 18968
rect 20710 18908 20736 18934
rect 24114 18942 24140 18968
rect 24436 18942 24462 18968
rect 23194 18908 23220 18934
rect 23240 18908 23266 18934
rect 24252 18908 24278 18934
rect 24344 18929 24370 18934
rect 24344 18912 24348 18929
rect 24348 18912 24365 18929
rect 24365 18912 24370 18929
rect 24344 18908 24370 18912
rect 25356 18929 25382 18934
rect 25356 18912 25360 18929
rect 25360 18912 25377 18929
rect 25377 18912 25382 18929
rect 25356 18908 25382 18912
rect 25494 18963 25520 18968
rect 25494 18946 25498 18963
rect 25498 18946 25515 18963
rect 25515 18946 25520 18963
rect 25494 18942 25520 18946
rect 26506 18963 26532 18968
rect 26506 18946 26508 18963
rect 26508 18946 26532 18963
rect 26506 18942 26532 18946
rect 25448 18929 25474 18934
rect 25448 18912 25452 18929
rect 25452 18912 25469 18929
rect 25469 18912 25474 18929
rect 25448 18908 25474 18912
rect 25632 18908 25658 18934
rect 25724 18908 25750 18934
rect 28024 18908 28050 18934
rect 28346 18929 28372 18934
rect 28346 18912 28367 18929
rect 28367 18912 28372 18929
rect 28346 18908 28372 18912
rect 28530 18908 28556 18934
rect 29588 18929 29614 18934
rect 29588 18912 29592 18929
rect 29592 18912 29609 18929
rect 29609 18912 29614 18929
rect 29588 18908 29614 18912
rect 29634 18929 29660 18934
rect 29634 18912 29638 18929
rect 29638 18912 29655 18929
rect 29655 18912 29660 18929
rect 29634 18908 29660 18912
rect 29680 18929 29706 18934
rect 29680 18912 29687 18929
rect 29687 18912 29704 18929
rect 29704 18912 29706 18929
rect 29680 18908 29706 18912
rect 4978 18806 5004 18832
rect 8566 18806 8592 18832
rect 9072 18806 9098 18832
rect 9532 18806 9558 18832
rect 13074 18806 13100 18832
rect 15696 18806 15722 18832
rect 19146 18806 19172 18832
rect 22918 18806 22944 18832
rect 24022 18840 24048 18866
rect 24298 18806 24324 18832
rect 24666 18806 24692 18832
rect 25494 18840 25520 18866
rect 29542 18895 29568 18900
rect 29542 18878 29546 18895
rect 29546 18878 29563 18895
rect 29563 18878 29568 18895
rect 29542 18874 29568 18878
rect 27978 18840 28004 18866
rect 27380 18806 27406 18832
rect 4840 18704 4866 18730
rect 5070 18602 5096 18628
rect 5668 18704 5694 18730
rect 10360 18704 10386 18730
rect 15742 18704 15768 18730
rect 12982 18670 13008 18696
rect 13672 18636 13698 18662
rect 5806 18602 5832 18628
rect 8290 18623 8316 18628
rect 8290 18606 8294 18623
rect 8294 18606 8311 18623
rect 8311 18606 8316 18623
rect 8290 18602 8316 18606
rect 8566 18602 8592 18628
rect 4656 18589 4682 18594
rect 4656 18572 4660 18589
rect 4660 18572 4677 18589
rect 4677 18572 4682 18589
rect 4656 18568 4682 18572
rect 4794 18589 4820 18594
rect 4794 18572 4798 18589
rect 4798 18572 4815 18589
rect 4815 18572 4820 18589
rect 4794 18568 4820 18572
rect 5484 18589 5510 18594
rect 5484 18572 5486 18589
rect 5486 18572 5510 18589
rect 5484 18568 5510 18572
rect 8520 18589 8546 18594
rect 8520 18572 8522 18589
rect 8522 18572 8546 18589
rect 9348 18602 9374 18628
rect 10774 18602 10800 18628
rect 11050 18623 11076 18628
rect 11050 18606 11057 18623
rect 11057 18606 11074 18623
rect 11074 18606 11076 18623
rect 11050 18602 11076 18606
rect 8520 18568 8546 18572
rect 10866 18589 10892 18594
rect 10866 18572 10870 18589
rect 10870 18572 10887 18589
rect 10887 18572 10892 18589
rect 10866 18568 10892 18572
rect 11004 18589 11030 18594
rect 11004 18572 11008 18589
rect 11008 18572 11025 18589
rect 11025 18572 11030 18589
rect 11004 18568 11030 18572
rect 5116 18534 5142 18560
rect 5254 18534 5280 18560
rect 6266 18534 6292 18560
rect 9486 18534 9512 18560
rect 10912 18534 10938 18560
rect 11832 18602 11858 18628
rect 13074 18623 13100 18628
rect 13074 18606 13078 18623
rect 13078 18606 13095 18623
rect 13095 18606 13100 18623
rect 13074 18602 13100 18606
rect 13120 18623 13146 18628
rect 13120 18606 13127 18623
rect 13127 18606 13144 18623
rect 13144 18606 13146 18623
rect 13120 18602 13146 18606
rect 13856 18602 13882 18628
rect 14086 18602 14112 18628
rect 15144 18636 15170 18662
rect 14316 18623 14342 18628
rect 14316 18606 14337 18623
rect 14337 18606 14342 18623
rect 14316 18602 14342 18606
rect 15052 18602 15078 18628
rect 15650 18636 15676 18662
rect 15788 18636 15814 18662
rect 15696 18623 15722 18628
rect 15696 18606 15700 18623
rect 15700 18606 15717 18623
rect 15717 18606 15722 18623
rect 15696 18602 15722 18606
rect 11464 18568 11490 18594
rect 11648 18589 11674 18594
rect 11648 18572 11650 18589
rect 11650 18572 11674 18589
rect 11648 18568 11674 18572
rect 14454 18568 14480 18594
rect 15236 18568 15262 18594
rect 18456 18636 18482 18662
rect 15972 18602 15998 18628
rect 16156 18623 16182 18628
rect 16156 18606 16160 18623
rect 16160 18606 16177 18623
rect 16177 18606 16182 18623
rect 16156 18602 16182 18606
rect 16202 18602 16228 18628
rect 19238 18623 19264 18628
rect 19238 18606 19242 18623
rect 19242 18606 19259 18623
rect 19259 18606 19264 18623
rect 19238 18602 19264 18606
rect 20664 18636 20690 18662
rect 19376 18623 19402 18628
rect 19376 18606 19397 18623
rect 19397 18606 19402 18623
rect 19376 18602 19402 18606
rect 20480 18602 20506 18628
rect 20618 18589 20644 18594
rect 20618 18572 20622 18589
rect 20622 18572 20639 18589
rect 20639 18572 20644 18589
rect 20618 18568 20644 18572
rect 20664 18589 20690 18594
rect 20664 18572 20668 18589
rect 20668 18572 20685 18589
rect 20685 18572 20690 18589
rect 20664 18568 20690 18572
rect 20940 18568 20966 18594
rect 13994 18534 14020 18560
rect 15742 18555 15768 18560
rect 15742 18538 15746 18555
rect 15746 18538 15763 18555
rect 15763 18538 15768 18555
rect 15742 18534 15768 18538
rect 15788 18555 15814 18560
rect 15788 18538 15792 18555
rect 15792 18538 15809 18555
rect 15809 18538 15814 18555
rect 15788 18534 15814 18538
rect 15834 18555 15860 18560
rect 15834 18538 15838 18555
rect 15838 18538 15855 18555
rect 15855 18538 15860 18555
rect 15834 18534 15860 18538
rect 17168 18534 17194 18560
rect 21262 18555 21288 18560
rect 21262 18538 21266 18555
rect 21266 18538 21283 18555
rect 21283 18538 21288 18555
rect 21262 18534 21288 18538
rect 22596 18704 22622 18730
rect 21952 18623 21978 18628
rect 21952 18606 21956 18623
rect 21956 18606 21973 18623
rect 21973 18606 21978 18623
rect 21952 18602 21978 18606
rect 22090 18623 22116 18628
rect 22826 18670 22852 18696
rect 25356 18704 25382 18730
rect 27288 18704 27314 18730
rect 25448 18670 25474 18696
rect 27058 18670 27084 18696
rect 22090 18606 22114 18623
rect 22114 18606 22116 18623
rect 22090 18602 22116 18606
rect 22366 18636 22392 18662
rect 24114 18636 24140 18662
rect 26230 18636 26256 18662
rect 22320 18602 22346 18628
rect 21354 18555 21380 18560
rect 21354 18538 21358 18555
rect 21358 18538 21375 18555
rect 21375 18538 21380 18555
rect 21354 18534 21380 18538
rect 23148 18568 23174 18594
rect 24160 18602 24186 18628
rect 24482 18589 24508 18594
rect 24482 18572 24484 18589
rect 24484 18572 24508 18589
rect 24482 18568 24508 18572
rect 26690 18602 26716 18628
rect 27978 18657 28004 18662
rect 27978 18640 27982 18657
rect 27982 18640 27999 18657
rect 27999 18640 28004 18657
rect 27978 18636 28004 18640
rect 27564 18623 27590 18628
rect 27564 18606 27571 18623
rect 27571 18606 27588 18623
rect 27588 18606 27590 18623
rect 27564 18602 27590 18606
rect 28300 18602 28326 18628
rect 26230 18589 26256 18594
rect 26230 18572 26234 18589
rect 26234 18572 26251 18589
rect 26251 18572 26256 18589
rect 26230 18568 26256 18572
rect 26276 18589 26302 18594
rect 26276 18572 26280 18589
rect 26280 18572 26297 18589
rect 26297 18572 26302 18589
rect 26276 18568 26302 18572
rect 27380 18589 27406 18594
rect 27380 18572 27384 18589
rect 27384 18572 27401 18589
rect 27401 18572 27406 18589
rect 27380 18568 27406 18572
rect 27518 18589 27544 18594
rect 27518 18572 27522 18589
rect 27522 18572 27539 18589
rect 27539 18572 27544 18589
rect 27518 18568 27544 18572
rect 28254 18568 28280 18594
rect 26460 18534 26486 18560
rect 28438 18534 28464 18560
rect 4794 18432 4820 18458
rect 4840 18432 4866 18458
rect 6036 18432 6062 18458
rect 6266 18453 6292 18458
rect 6266 18436 6270 18453
rect 6270 18436 6287 18453
rect 6287 18436 6292 18453
rect 6266 18432 6292 18436
rect 9532 18432 9558 18458
rect 3552 18419 3578 18424
rect 3552 18402 3554 18419
rect 3554 18402 3578 18419
rect 3552 18398 3578 18402
rect 11004 18432 11030 18458
rect 11648 18432 11674 18458
rect 12844 18432 12870 18458
rect 13994 18432 14020 18458
rect 14454 18432 14480 18458
rect 15788 18432 15814 18458
rect 17168 18432 17194 18458
rect 20664 18432 20690 18458
rect 21952 18432 21978 18458
rect 10222 18419 10248 18424
rect 3138 18364 3164 18390
rect 3598 18364 3624 18390
rect 5576 18364 5602 18390
rect 6174 18364 6200 18390
rect 6956 18364 6982 18390
rect 7002 18364 7028 18390
rect 7094 18364 7120 18390
rect 9302 18364 9328 18390
rect 9394 18385 9420 18390
rect 9394 18368 9409 18385
rect 9409 18368 9420 18385
rect 9394 18364 9420 18368
rect 9486 18385 9512 18390
rect 9486 18368 9503 18385
rect 9503 18368 9512 18385
rect 9547 18396 9573 18400
rect 9547 18379 9551 18396
rect 9551 18379 9568 18396
rect 9568 18379 9573 18396
rect 9547 18374 9573 18379
rect 9486 18364 9512 18368
rect 10222 18402 10224 18419
rect 10224 18402 10248 18419
rect 10222 18398 10248 18402
rect 12798 18398 12824 18424
rect 15052 18398 15078 18424
rect 5392 18330 5418 18356
rect 5300 18262 5326 18288
rect 9440 18296 9466 18322
rect 9486 18296 9512 18322
rect 6956 18262 6982 18288
rect 7278 18262 7304 18288
rect 7508 18262 7534 18288
rect 9210 18262 9236 18288
rect 10314 18364 10340 18390
rect 13074 18364 13100 18390
rect 13672 18364 13698 18390
rect 15236 18364 15262 18390
rect 15512 18364 15538 18390
rect 15742 18364 15768 18390
rect 12752 18330 12778 18356
rect 14454 18330 14480 18356
rect 15190 18351 15216 18356
rect 15190 18334 15194 18351
rect 15194 18334 15211 18351
rect 15211 18334 15216 18351
rect 15190 18330 15216 18334
rect 16524 18364 16550 18390
rect 17122 18364 17148 18390
rect 17214 18385 17240 18390
rect 17214 18368 17218 18385
rect 17218 18368 17235 18385
rect 17235 18368 17240 18385
rect 17214 18364 17240 18368
rect 17260 18385 17286 18390
rect 17260 18368 17267 18385
rect 17267 18368 17284 18385
rect 17284 18368 17286 18385
rect 17260 18364 17286 18368
rect 17950 18364 17976 18390
rect 18456 18385 18482 18390
rect 18456 18368 18477 18385
rect 18477 18368 18482 18385
rect 23056 18398 23082 18424
rect 24298 18419 24324 18424
rect 24298 18402 24302 18419
rect 24302 18402 24319 18419
rect 24319 18402 24324 18419
rect 24298 18398 24324 18402
rect 27518 18432 27544 18458
rect 28438 18432 28464 18458
rect 29634 18432 29660 18458
rect 28346 18398 28372 18424
rect 28622 18419 28648 18424
rect 28622 18402 28624 18419
rect 28624 18402 28648 18419
rect 28622 18398 28648 18402
rect 18456 18364 18482 18368
rect 18916 18364 18942 18390
rect 20664 18364 20690 18390
rect 21308 18364 21334 18390
rect 21630 18364 21656 18390
rect 22780 18364 22806 18390
rect 23148 18385 23174 18390
rect 23148 18368 23169 18385
rect 23169 18368 23174 18385
rect 23148 18364 23174 18368
rect 24390 18385 24416 18390
rect 24390 18368 24394 18385
rect 24394 18368 24411 18385
rect 24411 18368 24416 18385
rect 24390 18364 24416 18368
rect 24482 18385 24508 18390
rect 24482 18368 24489 18385
rect 24489 18368 24506 18385
rect 24506 18368 24508 18385
rect 24482 18364 24508 18368
rect 27564 18364 27590 18390
rect 29772 18364 29798 18390
rect 10176 18262 10202 18288
rect 14684 18262 14710 18288
rect 19238 18262 19264 18288
rect 22964 18330 22990 18356
rect 21078 18262 21104 18288
rect 24344 18351 24370 18356
rect 24344 18334 24348 18351
rect 24348 18334 24365 18351
rect 24365 18334 24370 18351
rect 24344 18330 24370 18334
rect 27978 18330 28004 18356
rect 24482 18296 24508 18322
rect 23148 18262 23174 18288
rect 24160 18262 24186 18288
rect 3598 18160 3624 18186
rect 4656 18160 4682 18186
rect 3138 18079 3164 18084
rect 3138 18062 3142 18079
rect 3142 18062 3159 18079
rect 3159 18062 3164 18079
rect 3138 18058 3164 18062
rect 5668 18160 5694 18186
rect 6036 18181 6062 18186
rect 6036 18164 6040 18181
rect 6040 18164 6057 18181
rect 6057 18164 6062 18181
rect 6036 18160 6062 18164
rect 6910 18160 6936 18186
rect 6772 18126 6798 18152
rect 9118 18160 9144 18186
rect 9486 18160 9512 18186
rect 10774 18160 10800 18186
rect 10866 18160 10892 18186
rect 5300 18113 5326 18118
rect 5300 18096 5304 18113
rect 5304 18096 5321 18113
rect 5321 18096 5326 18113
rect 5300 18092 5326 18096
rect 7554 18092 7580 18118
rect 3736 18058 3762 18084
rect 6680 18079 6706 18084
rect 6680 18062 6684 18079
rect 6684 18062 6701 18079
rect 6701 18062 6706 18079
rect 6680 18058 6706 18062
rect 6726 18058 6752 18084
rect 6864 18079 6890 18084
rect 6864 18062 6868 18079
rect 6868 18062 6885 18079
rect 6885 18062 6890 18079
rect 6864 18058 6890 18062
rect 5576 18024 5602 18050
rect 5990 18024 6016 18050
rect 6772 18045 6798 18050
rect 6772 18028 6776 18045
rect 6776 18028 6793 18045
rect 6793 18028 6798 18045
rect 6772 18024 6798 18028
rect 6818 18045 6844 18050
rect 6818 18028 6822 18045
rect 6822 18028 6839 18045
rect 6839 18028 6844 18045
rect 6818 18024 6844 18028
rect 7508 18058 7534 18084
rect 7646 18079 7672 18084
rect 7646 18062 7650 18079
rect 7650 18062 7667 18079
rect 7667 18062 7672 18079
rect 7646 18058 7672 18062
rect 7600 18045 7626 18050
rect 7600 18028 7604 18045
rect 7604 18028 7621 18045
rect 7621 18028 7626 18045
rect 7600 18024 7626 18028
rect 8290 18058 8316 18084
rect 8428 18079 8454 18084
rect 8428 18062 8432 18079
rect 8432 18062 8449 18079
rect 8449 18062 8454 18079
rect 8428 18058 8454 18062
rect 8566 18079 8592 18084
rect 8566 18062 8587 18079
rect 8587 18062 8592 18079
rect 8566 18058 8592 18062
rect 10176 18079 10202 18084
rect 10176 18062 10180 18079
rect 10180 18062 10197 18079
rect 10197 18062 10202 18079
rect 10176 18058 10202 18062
rect 10314 18079 10340 18084
rect 10314 18062 10335 18079
rect 10335 18062 10340 18079
rect 10314 18058 10340 18062
rect 12752 18058 12778 18084
rect 13856 18160 13882 18186
rect 14454 18160 14480 18186
rect 14684 18160 14710 18186
rect 14868 18126 14894 18152
rect 8336 18024 8362 18050
rect 10406 18045 10432 18050
rect 10406 18028 10408 18045
rect 10408 18028 10432 18045
rect 10406 18024 10432 18028
rect 12936 18024 12962 18050
rect 13074 18024 13100 18050
rect 13948 18058 13974 18084
rect 14684 18079 14710 18084
rect 14684 18062 14688 18079
rect 14688 18062 14705 18079
rect 14705 18062 14710 18079
rect 14684 18058 14710 18062
rect 14776 18079 14802 18084
rect 14776 18062 14782 18079
rect 14782 18062 14802 18079
rect 14776 18058 14802 18062
rect 17214 18160 17240 18186
rect 20526 18160 20552 18186
rect 15190 18092 15216 18118
rect 21124 18160 21150 18186
rect 21354 18160 21380 18186
rect 21446 18160 21472 18186
rect 21584 18160 21610 18186
rect 22090 18160 22116 18186
rect 23056 18160 23082 18186
rect 28300 18160 28326 18186
rect 28438 18160 28464 18186
rect 22320 18126 22346 18152
rect 27104 18126 27130 18152
rect 15006 18079 15032 18084
rect 15006 18062 15017 18079
rect 15017 18062 15032 18079
rect 15006 18058 15032 18062
rect 15052 18058 15078 18084
rect 16156 18058 16182 18084
rect 17720 18058 17746 18084
rect 20664 18058 20690 18084
rect 21078 18058 21104 18084
rect 23240 18092 23266 18118
rect 23424 18092 23450 18118
rect 21630 18058 21656 18084
rect 13626 18045 13652 18050
rect 13626 18028 13628 18045
rect 13628 18028 13652 18045
rect 13626 18024 13652 18028
rect 16478 18024 16504 18050
rect 21446 18045 21472 18050
rect 21446 18028 21448 18045
rect 21448 18028 21472 18045
rect 21446 18024 21472 18028
rect 7692 17990 7718 18016
rect 15052 17990 15078 18016
rect 19376 17990 19402 18016
rect 20158 17990 20184 18016
rect 14684 17888 14710 17914
rect 22366 17888 22392 17914
rect 24252 17909 24278 17914
rect 24252 17892 24256 17909
rect 24256 17892 24273 17909
rect 24273 17892 24278 17909
rect 24252 17888 24278 17892
rect 5760 17854 5786 17880
rect 6174 17854 6200 17880
rect 12430 17854 12456 17880
rect 13074 17854 13100 17880
rect 21354 17854 21380 17880
rect 22964 17875 22990 17880
rect 22964 17858 22966 17875
rect 22966 17858 22990 17875
rect 22964 17854 22990 17858
rect 26460 17875 26486 17880
rect 26460 17858 26462 17875
rect 26462 17858 26486 17875
rect 26460 17854 26486 17858
rect 6956 17820 6982 17846
rect 7002 17820 7028 17846
rect 12752 17820 12778 17846
rect 12936 17841 12962 17846
rect 12936 17824 12957 17841
rect 12957 17824 12962 17841
rect 12936 17820 12962 17824
rect 18778 17841 18804 17846
rect 18778 17824 18782 17841
rect 18782 17824 18799 17841
rect 18799 17824 18804 17841
rect 18778 17820 18804 17824
rect 18870 17841 18896 17846
rect 18870 17824 18874 17841
rect 18874 17824 18891 17841
rect 18891 17824 18896 17841
rect 18870 17820 18896 17824
rect 20158 17820 20184 17846
rect 20664 17820 20690 17846
rect 21492 17820 21518 17846
rect 22780 17820 22806 17846
rect 23976 17820 24002 17846
rect 24068 17841 24094 17846
rect 24068 17824 24083 17841
rect 24083 17824 24094 17841
rect 24068 17820 24094 17824
rect 7600 17786 7626 17812
rect 21078 17807 21104 17812
rect 21078 17790 21082 17807
rect 21082 17790 21099 17807
rect 21099 17790 21104 17807
rect 21078 17786 21104 17790
rect 19284 17718 19310 17744
rect 21216 17718 21242 17744
rect 21354 17718 21380 17744
rect 22458 17718 22484 17744
rect 23148 17718 23174 17744
rect 26138 17820 26164 17846
rect 26368 17841 26394 17846
rect 26368 17824 26389 17841
rect 26389 17824 26394 17841
rect 26368 17820 26394 17824
rect 26184 17786 26210 17812
rect 27104 17786 27130 17812
rect 27426 17786 27452 17812
rect 24298 17752 24324 17778
rect 25724 17718 25750 17744
rect 29588 17752 29614 17778
rect 27104 17718 27130 17744
rect 4702 17616 4728 17642
rect 6818 17616 6844 17642
rect 3138 17569 3164 17574
rect 3138 17552 3142 17569
rect 3142 17552 3159 17569
rect 3159 17552 3164 17569
rect 3138 17548 3164 17552
rect 8428 17616 8454 17642
rect 9394 17616 9420 17642
rect 18778 17637 18804 17642
rect 18778 17620 18782 17637
rect 18782 17620 18799 17637
rect 18799 17620 18804 17637
rect 18778 17616 18804 17620
rect 19008 17582 19034 17608
rect 20112 17582 20138 17608
rect 3184 17514 3210 17540
rect 4748 17535 4774 17540
rect 4748 17518 4752 17535
rect 4752 17518 4769 17535
rect 4769 17518 4774 17535
rect 4748 17514 4774 17518
rect 5208 17514 5234 17540
rect 5668 17514 5694 17540
rect 5760 17535 5786 17540
rect 5760 17518 5781 17535
rect 5781 17518 5786 17535
rect 5760 17514 5786 17518
rect 8566 17514 8592 17540
rect 3414 17480 3440 17506
rect 4794 17501 4820 17506
rect 4794 17484 4798 17501
rect 4798 17484 4815 17501
rect 4815 17484 4820 17501
rect 4794 17480 4820 17484
rect 5852 17501 5878 17506
rect 5852 17484 5854 17501
rect 5854 17484 5878 17501
rect 5852 17480 5878 17484
rect 8474 17501 8500 17506
rect 8474 17484 8476 17501
rect 8476 17484 8500 17501
rect 8474 17480 8500 17484
rect 11188 17446 11214 17472
rect 13902 17446 13928 17472
rect 14454 17446 14480 17472
rect 16202 17446 16228 17472
rect 18824 17535 18850 17540
rect 18824 17518 18839 17535
rect 18839 17518 18850 17535
rect 18824 17514 18850 17518
rect 18916 17535 18942 17540
rect 19146 17548 19172 17574
rect 18916 17518 18933 17535
rect 18933 17518 18942 17535
rect 18916 17514 18942 17518
rect 18991 17525 19017 17529
rect 18991 17508 18995 17525
rect 18995 17508 19012 17525
rect 19012 17508 19017 17525
rect 18991 17503 19017 17508
rect 19928 17514 19954 17540
rect 22918 17616 22944 17642
rect 24068 17616 24094 17642
rect 23976 17582 24002 17608
rect 21078 17548 21104 17574
rect 21216 17548 21242 17574
rect 22458 17569 22484 17574
rect 22458 17552 22462 17569
rect 22462 17552 22479 17569
rect 22479 17552 22484 17569
rect 22458 17548 22484 17552
rect 27242 17616 27268 17642
rect 26138 17582 26164 17608
rect 26322 17582 26348 17608
rect 26920 17582 26946 17608
rect 22780 17514 22806 17540
rect 23102 17514 23128 17540
rect 24160 17514 24186 17540
rect 24436 17514 24462 17540
rect 24620 17514 24646 17540
rect 25632 17514 25658 17540
rect 25770 17535 25796 17540
rect 25770 17518 25774 17535
rect 25774 17518 25791 17535
rect 25791 17518 25796 17535
rect 25770 17514 25796 17518
rect 19100 17446 19126 17472
rect 21630 17480 21656 17506
rect 22044 17480 22070 17506
rect 22688 17501 22714 17506
rect 22688 17484 22690 17501
rect 22690 17484 22714 17501
rect 22688 17480 22714 17484
rect 24528 17480 24554 17506
rect 26092 17535 26118 17540
rect 26092 17518 26103 17535
rect 26103 17518 26118 17535
rect 25862 17446 25888 17472
rect 26092 17514 26118 17518
rect 26184 17514 26210 17540
rect 26736 17514 26762 17540
rect 27978 17535 28004 17540
rect 27978 17518 27982 17535
rect 27982 17518 27999 17535
rect 27999 17518 28004 17535
rect 27978 17514 28004 17518
rect 29588 17514 29614 17540
rect 26368 17480 26394 17506
rect 28024 17480 28050 17506
rect 28208 17501 28234 17506
rect 28208 17484 28210 17501
rect 28210 17484 28234 17501
rect 28208 17480 28234 17484
rect 29496 17446 29522 17472
rect 4794 17344 4820 17370
rect 18916 17344 18942 17370
rect 26368 17344 26394 17370
rect 27334 17344 27360 17370
rect 3828 17331 3854 17336
rect 3828 17314 3830 17331
rect 3830 17314 3854 17331
rect 3828 17310 3854 17314
rect 7462 17331 7488 17336
rect 7462 17314 7464 17331
rect 7464 17314 7488 17331
rect 7462 17310 7488 17314
rect 12614 17310 12640 17336
rect 12844 17331 12870 17336
rect 12844 17314 12846 17331
rect 12846 17314 12870 17331
rect 12844 17310 12870 17314
rect 14454 17310 14480 17336
rect 17996 17310 18022 17336
rect 5760 17276 5786 17302
rect 6956 17276 6982 17302
rect 7232 17297 7258 17302
rect 7232 17280 7236 17297
rect 7236 17280 7253 17297
rect 7253 17280 7258 17297
rect 7232 17276 7258 17280
rect 7554 17276 7580 17302
rect 7876 17276 7902 17302
rect 12660 17276 12686 17302
rect 12936 17276 12962 17302
rect 13948 17276 13974 17302
rect 17720 17297 17746 17302
rect 17720 17280 17724 17297
rect 17724 17280 17741 17297
rect 17741 17280 17746 17297
rect 17720 17276 17746 17280
rect 17858 17297 17884 17302
rect 17858 17280 17879 17297
rect 17879 17280 17884 17297
rect 17858 17276 17884 17280
rect 19652 17276 19678 17302
rect 20158 17276 20184 17302
rect 23240 17310 23266 17336
rect 25586 17331 25612 17336
rect 25586 17314 25588 17331
rect 25588 17314 25612 17331
rect 25586 17310 25612 17314
rect 27058 17310 27084 17336
rect 20802 17276 20828 17302
rect 23102 17297 23128 17302
rect 23102 17280 23123 17297
rect 23123 17280 23128 17297
rect 23102 17276 23128 17280
rect 25632 17276 25658 17302
rect 27104 17297 27130 17302
rect 27104 17280 27108 17297
rect 27108 17280 27125 17297
rect 27125 17280 27130 17297
rect 27104 17276 27130 17280
rect 28438 17331 28464 17336
rect 28438 17314 28440 17331
rect 28440 17314 28464 17331
rect 28438 17310 28464 17314
rect 29496 17331 29522 17336
rect 29496 17314 29500 17331
rect 29500 17314 29517 17331
rect 29517 17314 29522 17331
rect 29496 17310 29522 17314
rect 27242 17297 27268 17302
rect 27242 17280 27266 17297
rect 27266 17280 27268 17297
rect 27242 17276 27268 17280
rect 27426 17297 27452 17302
rect 27426 17280 27437 17297
rect 27437 17280 27452 17297
rect 3138 17242 3164 17268
rect 8428 17208 8454 17234
rect 8658 17208 8684 17234
rect 10038 17208 10064 17234
rect 10176 17208 10202 17234
rect 10590 17208 10616 17234
rect 10912 17208 10938 17234
rect 14500 17242 14526 17268
rect 17030 17242 17056 17268
rect 17674 17242 17700 17268
rect 8290 17174 8316 17200
rect 9624 17174 9650 17200
rect 11648 17174 11674 17200
rect 14316 17174 14342 17200
rect 15236 17174 15262 17200
rect 20572 17174 20598 17200
rect 21446 17174 21472 17200
rect 24712 17242 24738 17268
rect 27426 17276 27452 17280
rect 24298 17208 24324 17234
rect 23148 17174 23174 17200
rect 27748 17242 27774 17268
rect 26782 17208 26808 17234
rect 28024 17276 28050 17302
rect 28346 17297 28372 17302
rect 28346 17280 28367 17297
rect 28367 17280 28372 17297
rect 28346 17276 28372 17280
rect 29404 17276 29430 17302
rect 27978 17242 28004 17268
rect 29772 17276 29798 17302
rect 26736 17174 26762 17200
rect 28622 17174 28648 17200
rect 29496 17195 29522 17200
rect 29496 17178 29500 17195
rect 29500 17178 29517 17195
rect 29517 17178 29522 17195
rect 29496 17174 29522 17178
rect 5668 17072 5694 17098
rect 6680 17072 6706 17098
rect 8658 17025 8684 17030
rect 8658 17008 8662 17025
rect 8662 17008 8679 17025
rect 8679 17008 8684 17025
rect 8658 17004 8684 17008
rect 5760 16970 5786 16996
rect 6082 16970 6108 16996
rect 7048 16970 7074 16996
rect 8980 16970 9006 16996
rect 11970 17072 11996 17098
rect 24436 17072 24462 17098
rect 10912 17004 10938 17030
rect 12246 16991 12272 16996
rect 12246 16974 12250 16991
rect 12250 16974 12267 16991
rect 12267 16974 12272 16991
rect 12246 16970 12272 16974
rect 12752 17004 12778 17030
rect 15006 17004 15032 17030
rect 21216 17025 21242 17030
rect 14730 16991 14756 16996
rect 14730 16974 14734 16991
rect 14734 16974 14751 16991
rect 14751 16974 14756 16991
rect 14730 16970 14756 16974
rect 7140 16936 7166 16962
rect 7462 16936 7488 16962
rect 8934 16936 8960 16962
rect 10130 16936 10156 16962
rect 10636 16936 10662 16962
rect 11188 16957 11214 16962
rect 11188 16940 11190 16957
rect 11190 16940 11214 16957
rect 11188 16936 11214 16940
rect 12936 16936 12962 16962
rect 13166 16957 13192 16962
rect 13166 16940 13168 16957
rect 13168 16940 13192 16957
rect 13166 16936 13192 16940
rect 14040 16936 14066 16962
rect 14776 16957 14802 16962
rect 14776 16940 14780 16957
rect 14780 16940 14797 16957
rect 14797 16940 14802 16957
rect 14776 16936 14802 16940
rect 15144 16991 15170 16996
rect 15144 16974 15148 16991
rect 15148 16974 15165 16991
rect 15165 16974 15170 16991
rect 15144 16970 15170 16974
rect 15236 16991 15262 16996
rect 15236 16974 15240 16991
rect 15240 16974 15257 16991
rect 15257 16974 15262 16991
rect 15236 16970 15262 16974
rect 15466 16970 15492 16996
rect 17122 16970 17148 16996
rect 17168 16991 17194 16996
rect 17168 16974 17172 16991
rect 17172 16974 17189 16991
rect 17189 16974 17194 16991
rect 17168 16970 17194 16974
rect 20572 16970 20598 16996
rect 21216 17008 21220 17025
rect 21220 17008 21237 17025
rect 21237 17008 21242 17025
rect 21216 17004 21242 17008
rect 24712 17072 24738 17098
rect 25770 17072 25796 17098
rect 26138 17072 26164 17098
rect 26966 17072 26992 17098
rect 27748 17072 27774 17098
rect 27978 17072 28004 17098
rect 28392 17072 28418 17098
rect 21492 16970 21518 16996
rect 21538 16970 21564 16996
rect 24574 16970 24600 16996
rect 15650 16936 15676 16962
rect 15834 16936 15860 16962
rect 16018 16957 16044 16962
rect 16018 16940 16020 16957
rect 16020 16940 16044 16957
rect 16018 16936 16044 16940
rect 22688 16936 22714 16962
rect 26736 16991 26762 16996
rect 26736 16974 26740 16991
rect 26740 16974 26757 16991
rect 26757 16974 26762 16991
rect 26736 16970 26762 16974
rect 28622 17025 28648 17030
rect 28622 17008 28626 17025
rect 28626 17008 28643 17025
rect 28643 17008 28648 17025
rect 28622 17004 28648 17008
rect 28300 16970 28326 16996
rect 29496 16970 29522 16996
rect 26414 16936 26440 16962
rect 26782 16936 26808 16962
rect 26966 16957 26992 16962
rect 26966 16940 26968 16957
rect 26968 16940 26992 16957
rect 26966 16936 26992 16940
rect 9532 16902 9558 16928
rect 12108 16902 12134 16928
rect 14270 16902 14296 16928
rect 14868 16902 14894 16928
rect 17076 16902 17102 16928
rect 17306 16902 17332 16928
rect 21676 16902 21702 16928
rect 28116 16902 28142 16928
rect 28990 16957 29016 16962
rect 28990 16940 28994 16957
rect 28994 16940 29011 16957
rect 29011 16940 29016 16957
rect 28990 16936 29016 16940
rect 29496 16902 29522 16928
rect 14040 16800 14066 16826
rect 15006 16821 15032 16826
rect 15006 16804 15010 16821
rect 15010 16804 15027 16821
rect 15027 16804 15032 16821
rect 15006 16800 15032 16804
rect 15052 16821 15078 16826
rect 15052 16804 15056 16821
rect 15056 16804 15073 16821
rect 15073 16804 15078 16821
rect 15052 16800 15078 16804
rect 18824 16800 18850 16826
rect 21262 16800 21288 16826
rect 22688 16800 22714 16826
rect 23010 16800 23036 16826
rect 27242 16800 27268 16826
rect 7554 16732 7580 16758
rect 8934 16766 8960 16792
rect 11648 16787 11674 16792
rect 11648 16770 11652 16787
rect 11652 16770 11669 16787
rect 11669 16770 11674 16787
rect 11648 16766 11674 16770
rect 12292 16766 12318 16792
rect 12660 16766 12686 16792
rect 13028 16787 13054 16792
rect 13028 16770 13030 16787
rect 13030 16770 13054 16787
rect 13028 16766 13054 16770
rect 14270 16766 14296 16792
rect 8336 16732 8362 16758
rect 8428 16732 8454 16758
rect 9532 16753 9558 16758
rect 9532 16736 9536 16753
rect 9536 16736 9553 16753
rect 9553 16736 9558 16753
rect 9532 16732 9558 16736
rect 9624 16753 9650 16758
rect 9624 16736 9628 16753
rect 9628 16736 9645 16753
rect 9645 16736 9650 16753
rect 9624 16732 9650 16736
rect 9670 16753 9696 16758
rect 9670 16736 9674 16753
rect 9674 16736 9691 16753
rect 9691 16736 9696 16753
rect 9670 16732 9696 16736
rect 7278 16719 7304 16724
rect 7278 16702 7282 16719
rect 7282 16702 7299 16719
rect 7299 16702 7304 16719
rect 7278 16698 7304 16702
rect 8382 16698 8408 16724
rect 10038 16753 10064 16758
rect 10038 16736 10042 16753
rect 10042 16736 10059 16753
rect 10059 16736 10064 16753
rect 10038 16732 10064 16736
rect 10176 16753 10202 16758
rect 10176 16736 10197 16753
rect 10197 16736 10202 16753
rect 10176 16732 10202 16736
rect 11694 16753 11720 16758
rect 11694 16736 11698 16753
rect 11698 16736 11715 16753
rect 11715 16736 11720 16753
rect 11694 16732 11720 16736
rect 11740 16753 11766 16758
rect 11740 16736 11747 16753
rect 11747 16736 11764 16753
rect 11764 16736 11766 16753
rect 11740 16732 11766 16736
rect 12108 16753 12134 16758
rect 12108 16736 12112 16753
rect 12112 16736 12129 16753
rect 12129 16736 12134 16753
rect 12108 16732 12134 16736
rect 12752 16732 12778 16758
rect 12844 16732 12870 16758
rect 12936 16753 12962 16758
rect 12936 16736 12957 16753
rect 12957 16736 12962 16753
rect 12936 16732 12962 16736
rect 14316 16753 14342 16758
rect 14316 16736 14320 16753
rect 14320 16736 14337 16753
rect 14337 16736 14342 16753
rect 14316 16732 14342 16736
rect 13856 16698 13882 16724
rect 14086 16698 14112 16724
rect 14454 16753 14480 16758
rect 14868 16787 14894 16792
rect 14868 16770 14872 16787
rect 14872 16770 14889 16787
rect 14889 16770 14894 16787
rect 14868 16766 14894 16770
rect 15558 16766 15584 16792
rect 17076 16787 17102 16792
rect 17076 16770 17080 16787
rect 17080 16770 17097 16787
rect 17097 16770 17102 16787
rect 17076 16766 17102 16770
rect 14454 16736 14471 16753
rect 14471 16736 14480 16753
rect 14454 16732 14480 16736
rect 14638 16753 14664 16758
rect 14638 16736 14649 16753
rect 14649 16736 14664 16753
rect 14638 16732 14664 16736
rect 15512 16732 15538 16758
rect 15834 16732 15860 16758
rect 15972 16732 15998 16758
rect 15190 16698 15216 16724
rect 15466 16698 15492 16724
rect 17122 16732 17148 16758
rect 17260 16766 17286 16792
rect 17720 16732 17746 16758
rect 17904 16732 17930 16758
rect 20112 16743 20138 16769
rect 20158 16753 20184 16758
rect 20158 16736 20179 16753
rect 20179 16736 20184 16753
rect 20158 16732 20184 16736
rect 20756 16732 20782 16758
rect 21308 16753 21334 16758
rect 21308 16736 21312 16753
rect 21312 16736 21329 16753
rect 21329 16736 21334 16753
rect 21308 16732 21334 16736
rect 4748 16630 4774 16656
rect 5024 16630 5050 16656
rect 6312 16630 6338 16656
rect 8382 16630 8408 16656
rect 9808 16651 9834 16656
rect 9808 16634 9812 16651
rect 9812 16634 9829 16651
rect 9829 16634 9834 16651
rect 9808 16630 9834 16634
rect 14546 16664 14572 16690
rect 16524 16664 16550 16690
rect 21446 16753 21472 16758
rect 21676 16766 21702 16792
rect 22918 16766 22944 16792
rect 26000 16766 26026 16792
rect 28346 16766 28372 16792
rect 28668 16766 28694 16792
rect 21446 16736 21463 16753
rect 21463 16736 21472 16753
rect 21446 16732 21472 16736
rect 22688 16732 22714 16758
rect 22780 16732 22806 16758
rect 23102 16753 23128 16758
rect 23102 16736 23123 16753
rect 23123 16736 23128 16753
rect 23102 16732 23128 16736
rect 26046 16732 26072 16758
rect 26414 16732 26440 16758
rect 28392 16753 28418 16758
rect 28392 16736 28396 16753
rect 28396 16736 28413 16753
rect 28413 16736 28418 16753
rect 28392 16732 28418 16736
rect 11740 16630 11766 16656
rect 12154 16630 12180 16656
rect 12798 16630 12824 16656
rect 13028 16630 13054 16656
rect 15880 16630 15906 16656
rect 17214 16630 17240 16656
rect 21906 16664 21932 16690
rect 20572 16630 20598 16656
rect 23148 16630 23174 16656
rect 24114 16630 24140 16656
rect 26690 16630 26716 16656
rect 29634 16630 29660 16656
rect 4748 16528 4774 16554
rect 4702 16494 4728 16520
rect 6772 16528 6798 16554
rect 9670 16528 9696 16554
rect 4656 16447 4682 16452
rect 4656 16430 4660 16447
rect 4660 16430 4677 16447
rect 4677 16430 4682 16447
rect 4656 16426 4682 16430
rect 4748 16447 4774 16452
rect 4748 16430 4754 16447
rect 4754 16430 4774 16447
rect 4748 16426 4774 16430
rect 3690 16392 3716 16418
rect 4564 16392 4590 16418
rect 4610 16392 4636 16418
rect 4917 16447 4943 16452
rect 4917 16430 4921 16447
rect 4921 16430 4938 16447
rect 4938 16430 4943 16447
rect 4917 16426 4943 16430
rect 5668 16426 5694 16452
rect 7278 16460 7304 16486
rect 9854 16494 9880 16520
rect 11694 16528 11720 16554
rect 12476 16528 12502 16554
rect 12246 16494 12272 16520
rect 6312 16426 6338 16452
rect 7232 16426 7258 16452
rect 7416 16447 7442 16452
rect 7416 16430 7420 16447
rect 7420 16430 7437 16447
rect 7437 16430 7442 16447
rect 7416 16426 7442 16430
rect 8612 16426 8638 16452
rect 5622 16392 5648 16418
rect 5990 16392 6016 16418
rect 7186 16392 7212 16418
rect 8934 16392 8960 16418
rect 9808 16426 9834 16452
rect 10590 16481 10616 16486
rect 10590 16464 10594 16481
rect 10594 16464 10611 16481
rect 10611 16464 10616 16481
rect 10590 16460 10616 16464
rect 12752 16460 12778 16486
rect 13166 16426 13192 16452
rect 13948 16447 13974 16452
rect 13948 16430 13969 16447
rect 13969 16430 13974 16447
rect 13948 16426 13974 16430
rect 14500 16426 14526 16452
rect 14776 16528 14802 16554
rect 17168 16528 17194 16554
rect 20802 16528 20828 16554
rect 22918 16528 22944 16554
rect 24022 16528 24048 16554
rect 29496 16549 29522 16554
rect 29496 16532 29500 16549
rect 29500 16532 29517 16549
rect 29517 16532 29522 16549
rect 29496 16528 29522 16532
rect 24712 16494 24738 16520
rect 25586 16494 25612 16520
rect 15466 16460 15492 16486
rect 16202 16426 16228 16452
rect 17214 16447 17240 16452
rect 17214 16430 17218 16447
rect 17218 16430 17235 16447
rect 17235 16430 17240 16447
rect 17214 16426 17240 16430
rect 17306 16447 17332 16452
rect 17306 16430 17310 16447
rect 17310 16430 17327 16447
rect 17327 16430 17332 16447
rect 17306 16426 17332 16430
rect 21308 16426 21334 16452
rect 15926 16392 15952 16418
rect 23976 16413 24002 16418
rect 23976 16396 23980 16413
rect 23980 16396 23997 16413
rect 23997 16396 24002 16413
rect 23976 16392 24002 16396
rect 24114 16447 24140 16452
rect 24114 16430 24118 16447
rect 24118 16430 24135 16447
rect 24135 16430 24140 16447
rect 24114 16426 24140 16430
rect 26092 16426 26118 16452
rect 29588 16447 29614 16452
rect 29588 16430 29592 16447
rect 29592 16430 29609 16447
rect 29609 16430 29614 16447
rect 29588 16426 29614 16430
rect 29634 16447 29660 16452
rect 29634 16430 29638 16447
rect 29638 16430 29655 16447
rect 29655 16430 29660 16447
rect 29634 16426 29660 16430
rect 29680 16447 29706 16452
rect 29680 16430 29687 16447
rect 29687 16430 29704 16447
rect 29704 16430 29706 16447
rect 29680 16426 29706 16430
rect 29818 16426 29844 16452
rect 25862 16392 25888 16418
rect 29496 16413 29522 16418
rect 29496 16396 29500 16413
rect 29500 16396 29517 16413
rect 29517 16396 29522 16413
rect 29496 16392 29522 16396
rect 6726 16358 6752 16384
rect 10268 16379 10294 16384
rect 10268 16362 10272 16379
rect 10272 16362 10289 16379
rect 10289 16362 10294 16379
rect 10268 16358 10294 16362
rect 10636 16358 10662 16384
rect 17260 16379 17286 16384
rect 17260 16362 17264 16379
rect 17264 16362 17281 16379
rect 17281 16362 17286 16379
rect 17260 16358 17286 16362
rect 4288 16256 4314 16282
rect 5024 16256 5050 16282
rect 4564 16222 4590 16248
rect 6726 16277 6752 16282
rect 6726 16260 6730 16277
rect 6730 16260 6747 16277
rect 6747 16260 6752 16277
rect 6726 16256 6752 16260
rect 10268 16256 10294 16282
rect 14454 16256 14480 16282
rect 23976 16256 24002 16282
rect 29496 16256 29522 16282
rect 9026 16243 9052 16248
rect 3138 16188 3164 16214
rect 3368 16209 3394 16214
rect 3368 16192 3389 16209
rect 3389 16192 3394 16209
rect 3368 16188 3394 16192
rect 4472 16188 4498 16214
rect 4518 16209 4544 16214
rect 4518 16192 4522 16209
rect 4522 16192 4539 16209
rect 4539 16192 4544 16209
rect 4518 16188 4544 16192
rect 4794 16188 4820 16214
rect 6266 16209 6292 16214
rect 6266 16192 6270 16209
rect 6270 16192 6287 16209
rect 6287 16192 6292 16209
rect 6266 16188 6292 16192
rect 6312 16209 6338 16214
rect 6312 16192 6316 16209
rect 6316 16192 6333 16209
rect 6333 16192 6338 16209
rect 6312 16188 6338 16192
rect 6772 16209 6798 16214
rect 6772 16192 6776 16209
rect 6776 16192 6793 16209
rect 6793 16192 6798 16209
rect 6772 16188 6798 16192
rect 7278 16188 7304 16214
rect 7508 16188 7534 16214
rect 9026 16226 9028 16243
rect 9028 16226 9052 16243
rect 9026 16222 9052 16226
rect 12936 16243 12962 16248
rect 12936 16226 12938 16243
rect 12938 16226 12962 16243
rect 12936 16222 12962 16226
rect 20802 16222 20828 16248
rect 8244 16188 8270 16214
rect 8474 16188 8500 16214
rect 8612 16188 8638 16214
rect 8934 16209 8960 16214
rect 8934 16192 8955 16209
rect 8955 16192 8960 16209
rect 8934 16188 8960 16192
rect 12752 16188 12778 16214
rect 12844 16209 12870 16214
rect 12844 16192 12865 16209
rect 12865 16192 12870 16209
rect 12844 16188 12870 16192
rect 21032 16188 21058 16214
rect 20572 16154 20598 16180
rect 7186 16120 7212 16146
rect 22780 16188 22806 16214
rect 25908 16222 25934 16248
rect 28300 16222 28326 16248
rect 24528 16188 24554 16214
rect 26046 16209 26072 16214
rect 26046 16192 26067 16209
rect 26067 16192 26072 16209
rect 26046 16188 26072 16192
rect 28346 16188 28372 16214
rect 4518 16086 4544 16112
rect 5392 16086 5418 16112
rect 6634 16107 6660 16112
rect 6634 16090 6638 16107
rect 6638 16090 6655 16107
rect 6655 16090 6660 16107
rect 6634 16086 6660 16090
rect 8198 16086 8224 16112
rect 20756 16086 20782 16112
rect 21860 16086 21886 16112
rect 25356 16154 25382 16180
rect 23148 16086 23174 16112
rect 28300 16175 28326 16180
rect 28300 16158 28304 16175
rect 28304 16158 28321 16175
rect 28321 16158 28326 16175
rect 28300 16154 28326 16158
rect 26736 16086 26762 16112
rect 27196 16086 27222 16112
rect 4656 15984 4682 16010
rect 6266 15984 6292 16010
rect 3138 15937 3164 15942
rect 3138 15920 3142 15937
rect 3142 15920 3159 15937
rect 3159 15920 3164 15937
rect 3138 15916 3164 15920
rect 3414 15882 3440 15908
rect 4794 15882 4820 15908
rect 5714 15882 5740 15908
rect 5760 15882 5786 15908
rect 7508 15882 7534 15908
rect 8980 15984 9006 16010
rect 9302 15984 9328 16010
rect 8290 15950 8316 15976
rect 25816 15950 25842 15976
rect 8198 15903 8224 15908
rect 8198 15886 8204 15903
rect 8204 15886 8224 15903
rect 8198 15882 8224 15886
rect 3368 15869 3394 15874
rect 3368 15852 3370 15869
rect 3370 15852 3394 15869
rect 3368 15848 3394 15852
rect 5208 15848 5234 15874
rect 5392 15869 5418 15874
rect 5392 15852 5394 15869
rect 5394 15852 5418 15869
rect 5392 15848 5418 15852
rect 9210 15882 9236 15908
rect 9348 15848 9374 15874
rect 10774 15903 10800 15908
rect 10774 15886 10778 15903
rect 10778 15886 10795 15903
rect 10795 15886 10800 15903
rect 10774 15882 10800 15886
rect 25356 15916 25382 15942
rect 25586 15916 25612 15942
rect 25862 15916 25888 15942
rect 24160 15882 24186 15908
rect 25632 15903 25658 15908
rect 25632 15886 25636 15903
rect 25636 15886 25653 15903
rect 25653 15886 25658 15903
rect 25632 15882 25658 15886
rect 25724 15903 25750 15908
rect 25724 15886 25730 15903
rect 25730 15886 25750 15903
rect 25724 15882 25750 15886
rect 26092 15916 26118 15942
rect 26736 15937 26762 15942
rect 26736 15920 26740 15937
rect 26740 15920 26757 15937
rect 26757 15920 26762 15937
rect 26736 15916 26762 15920
rect 10820 15848 10846 15874
rect 24390 15848 24416 15874
rect 24574 15869 24600 15874
rect 24574 15852 24576 15869
rect 24576 15852 24600 15869
rect 24574 15848 24600 15852
rect 26368 15882 26394 15908
rect 28162 15882 28188 15908
rect 29312 15916 29338 15942
rect 26046 15848 26072 15874
rect 26782 15848 26808 15874
rect 27012 15848 27038 15874
rect 7232 15814 7258 15840
rect 8244 15814 8270 15840
rect 8336 15814 8362 15840
rect 8382 15814 8408 15840
rect 10636 15814 10662 15840
rect 11832 15814 11858 15840
rect 20986 15814 21012 15840
rect 22964 15814 22990 15840
rect 26506 15814 26532 15840
rect 27288 15814 27314 15840
rect 28760 15869 28786 15874
rect 28760 15852 28764 15869
rect 28764 15852 28781 15869
rect 28781 15852 28786 15869
rect 28760 15848 28786 15852
rect 28990 15882 29016 15908
rect 4610 15712 4636 15738
rect 5208 15712 5234 15738
rect 5622 15712 5648 15738
rect 21860 15712 21886 15738
rect 26368 15712 26394 15738
rect 28162 15712 28188 15738
rect 3690 15699 3716 15704
rect 3690 15682 3692 15699
rect 3692 15682 3716 15699
rect 3690 15678 3716 15682
rect 8428 15678 8454 15704
rect 3414 15644 3440 15670
rect 5668 15644 5694 15670
rect 5760 15644 5786 15670
rect 9026 15644 9052 15670
rect 9256 15644 9282 15670
rect 11096 15678 11122 15704
rect 12522 15644 12548 15670
rect 15374 15678 15400 15704
rect 13028 15644 13054 15670
rect 15466 15665 15492 15670
rect 18594 15678 18620 15704
rect 20112 15678 20138 15704
rect 20296 15699 20322 15704
rect 20296 15682 20298 15699
rect 20298 15682 20322 15699
rect 20296 15678 20322 15682
rect 24390 15678 24416 15704
rect 25586 15699 25612 15704
rect 15466 15648 15487 15665
rect 15487 15648 15492 15665
rect 15466 15644 15492 15648
rect 16202 15644 16228 15670
rect 18732 15644 18758 15670
rect 20802 15644 20828 15670
rect 21630 15665 21656 15670
rect 21630 15648 21645 15665
rect 21645 15648 21656 15665
rect 21630 15644 21656 15648
rect 21722 15665 21748 15670
rect 21722 15648 21739 15665
rect 21739 15648 21748 15665
rect 21722 15644 21748 15648
rect 21906 15665 21932 15670
rect 21906 15648 21917 15665
rect 21917 15648 21932 15665
rect 3138 15610 3164 15636
rect 3460 15631 3486 15636
rect 3460 15614 3464 15631
rect 3464 15614 3481 15631
rect 3481 15614 3486 15631
rect 3460 15610 3486 15614
rect 9118 15610 9144 15636
rect 12384 15610 12410 15636
rect 15190 15610 15216 15636
rect 18318 15631 18344 15636
rect 18318 15614 18322 15631
rect 18322 15614 18339 15631
rect 18339 15614 18344 15631
rect 18318 15610 18344 15614
rect 10452 15542 10478 15568
rect 13672 15542 13698 15568
rect 16248 15542 16274 15568
rect 18318 15542 18344 15568
rect 19974 15542 20000 15568
rect 21032 15610 21058 15636
rect 21400 15610 21426 15636
rect 21906 15644 21932 15648
rect 25356 15665 25382 15670
rect 25356 15648 25360 15665
rect 25360 15648 25377 15665
rect 25377 15648 25382 15665
rect 25356 15644 25382 15648
rect 25586 15682 25588 15699
rect 25588 15682 25612 15699
rect 25586 15678 25612 15682
rect 26046 15644 26072 15670
rect 26920 15644 26946 15670
rect 27104 15644 27130 15670
rect 27196 15665 27222 15670
rect 27196 15648 27211 15665
rect 27211 15648 27222 15665
rect 27196 15644 27222 15648
rect 27288 15668 27314 15670
rect 27288 15651 27305 15668
rect 27305 15651 27314 15668
rect 27288 15644 27314 15651
rect 27349 15665 27375 15670
rect 27349 15648 27353 15665
rect 27353 15648 27370 15665
rect 27370 15648 27375 15665
rect 27349 15644 27375 15648
rect 27564 15644 27590 15670
rect 27748 15610 27774 15636
rect 26506 15576 26532 15602
rect 28116 15576 28142 15602
rect 20250 15542 20276 15568
rect 20296 15542 20322 15568
rect 20388 15542 20414 15568
rect 22826 15542 22852 15568
rect 26000 15542 26026 15568
rect 26322 15542 26348 15568
rect 27104 15542 27130 15568
rect 27334 15542 27360 15568
rect 5714 15440 5740 15466
rect 15926 15440 15952 15466
rect 16432 15440 16458 15466
rect 16938 15440 16964 15466
rect 10774 15372 10800 15398
rect 5622 15338 5648 15364
rect 5990 15338 6016 15364
rect 7278 15338 7304 15364
rect 7416 15338 7442 15364
rect 5852 15304 5878 15330
rect 7002 15304 7028 15330
rect 7094 15304 7120 15330
rect 7784 15304 7810 15330
rect 8106 15338 8132 15364
rect 8428 15338 8454 15364
rect 10912 15338 10938 15364
rect 11142 15338 11168 15364
rect 13258 15338 13284 15364
rect 13810 15359 13836 15364
rect 13810 15342 13814 15359
rect 13814 15342 13831 15359
rect 13831 15342 13836 15359
rect 13810 15338 13836 15342
rect 13948 15359 13974 15364
rect 16064 15372 16090 15398
rect 16156 15372 16182 15398
rect 18916 15440 18942 15466
rect 20066 15440 20092 15466
rect 22642 15440 22668 15466
rect 20204 15406 20230 15432
rect 25678 15440 25704 15466
rect 27748 15440 27774 15466
rect 18318 15372 18344 15398
rect 13948 15342 13969 15359
rect 13969 15342 13974 15359
rect 13948 15338 13974 15342
rect 15972 15359 15998 15364
rect 15972 15342 15979 15359
rect 15979 15342 15996 15359
rect 15996 15342 15998 15359
rect 15972 15338 15998 15342
rect 16110 15338 16136 15364
rect 16892 15338 16918 15364
rect 16938 15359 16964 15364
rect 16938 15342 16942 15359
rect 16942 15342 16959 15359
rect 16959 15342 16964 15359
rect 16938 15338 16964 15342
rect 18732 15338 18758 15364
rect 11096 15325 11122 15330
rect 11096 15308 11098 15325
rect 11098 15308 11122 15325
rect 11096 15304 11122 15308
rect 14040 15325 14066 15330
rect 14040 15308 14042 15325
rect 14042 15308 14066 15325
rect 14040 15304 14066 15308
rect 15788 15325 15814 15330
rect 15788 15308 15792 15325
rect 15792 15308 15809 15325
rect 15809 15308 15814 15325
rect 15788 15304 15814 15308
rect 16202 15304 16228 15330
rect 16248 15325 16274 15330
rect 16248 15308 16252 15325
rect 16252 15308 16269 15325
rect 16269 15308 16274 15325
rect 16248 15304 16274 15308
rect 16340 15325 16366 15330
rect 16340 15308 16344 15325
rect 16344 15308 16361 15325
rect 16361 15308 16366 15325
rect 16340 15304 16366 15308
rect 16386 15325 16412 15330
rect 16386 15308 16390 15325
rect 16390 15308 16407 15325
rect 16407 15308 16412 15325
rect 16386 15304 16412 15308
rect 16570 15304 16596 15330
rect 17168 15325 17194 15330
rect 17168 15308 17170 15325
rect 17170 15308 17194 15325
rect 17168 15304 17194 15308
rect 18686 15325 18712 15330
rect 18686 15308 18688 15325
rect 18688 15308 18712 15325
rect 18870 15338 18896 15364
rect 18686 15304 18712 15308
rect 19974 15325 20000 15330
rect 19974 15308 19978 15325
rect 19978 15308 19995 15325
rect 19995 15308 20000 15325
rect 19974 15304 20000 15308
rect 20066 15325 20092 15330
rect 20066 15308 20070 15325
rect 20070 15308 20087 15325
rect 20087 15308 20092 15325
rect 20066 15304 20092 15308
rect 20204 15304 20230 15330
rect 25724 15406 25750 15432
rect 22826 15393 22852 15398
rect 22826 15376 22830 15393
rect 22830 15376 22847 15393
rect 22847 15376 22852 15393
rect 22826 15372 22852 15376
rect 24160 15372 24186 15398
rect 26736 15393 26762 15398
rect 26736 15376 26740 15393
rect 26740 15376 26757 15393
rect 26757 15376 26762 15393
rect 26736 15372 26762 15376
rect 20940 15338 20966 15364
rect 22872 15338 22898 15364
rect 22918 15359 22944 15364
rect 22918 15342 22922 15359
rect 22922 15342 22939 15359
rect 22939 15342 22944 15359
rect 22918 15338 22944 15342
rect 24390 15359 24416 15364
rect 24390 15342 24411 15359
rect 24411 15342 24416 15359
rect 24390 15338 24416 15342
rect 26782 15338 26808 15364
rect 22964 15304 22990 15330
rect 26966 15325 26992 15330
rect 26966 15308 26968 15325
rect 26968 15308 26992 15325
rect 26966 15304 26992 15308
rect 6772 15270 6798 15296
rect 9072 15270 9098 15296
rect 11970 15270 11996 15296
rect 14822 15270 14848 15296
rect 22872 15291 22898 15296
rect 22872 15274 22876 15291
rect 22876 15274 22893 15291
rect 22893 15274 22898 15291
rect 22872 15270 22898 15274
rect 5944 15168 5970 15194
rect 3782 15155 3808 15160
rect 3782 15138 3784 15155
rect 3784 15138 3808 15155
rect 3782 15134 3808 15138
rect 5162 15134 5188 15160
rect 6864 15155 6890 15160
rect 6864 15138 6868 15155
rect 6868 15138 6885 15155
rect 6885 15138 6890 15155
rect 6864 15134 6890 15138
rect 7140 15168 7166 15194
rect 3414 15100 3440 15126
rect 4840 15121 4866 15126
rect 4840 15104 4844 15121
rect 4844 15104 4861 15121
rect 4861 15104 4866 15121
rect 4840 15100 4866 15104
rect 4978 15121 5004 15126
rect 4978 15104 4982 15121
rect 4982 15104 4999 15121
rect 4999 15104 5004 15121
rect 4978 15100 5004 15104
rect 5070 15100 5096 15126
rect 3460 15066 3486 15092
rect 6450 15100 6476 15126
rect 6634 15100 6660 15126
rect 6772 15121 6798 15126
rect 6772 15104 6776 15121
rect 6776 15104 6793 15121
rect 6793 15104 6798 15121
rect 6772 15100 6798 15104
rect 6910 15121 6936 15126
rect 6910 15104 6914 15121
rect 6914 15104 6931 15121
rect 6931 15104 6936 15121
rect 6910 15100 6936 15104
rect 7048 15134 7074 15160
rect 7324 15100 7350 15126
rect 8980 15168 9006 15194
rect 9072 15168 9098 15194
rect 10544 15168 10570 15194
rect 7830 15100 7856 15126
rect 8842 15121 8868 15126
rect 8842 15104 8857 15121
rect 8857 15104 8868 15121
rect 8842 15100 8868 15104
rect 7278 15087 7304 15092
rect 7278 15070 7282 15087
rect 7282 15070 7299 15087
rect 7299 15070 7304 15087
rect 7278 15066 7304 15070
rect 9210 15100 9236 15126
rect 9164 15066 9190 15092
rect 4702 15032 4728 15058
rect 5024 15032 5050 15058
rect 8888 15032 8914 15058
rect 10268 15134 10294 15160
rect 10912 15100 10938 15126
rect 4794 14998 4820 15024
rect 5116 15019 5142 15024
rect 5116 15002 5120 15019
rect 5120 15002 5137 15019
rect 5137 15002 5142 15019
rect 5116 14998 5142 15002
rect 6404 15019 6430 15024
rect 6404 15002 6408 15019
rect 6408 15002 6425 15019
rect 6425 15002 6430 15019
rect 6404 14998 6430 15002
rect 7416 14998 7442 15024
rect 7462 14998 7488 15024
rect 9118 14998 9144 15024
rect 11832 15121 11858 15126
rect 11970 15168 11996 15194
rect 16386 15168 16412 15194
rect 21722 15168 21748 15194
rect 12844 15134 12870 15160
rect 13028 15155 13054 15160
rect 13028 15138 13030 15155
rect 13030 15138 13054 15155
rect 13028 15134 13054 15138
rect 11832 15104 11849 15121
rect 11849 15104 11858 15121
rect 11832 15100 11858 15104
rect 12062 15100 12088 15126
rect 12108 15066 12134 15092
rect 12384 15066 12410 15092
rect 13718 15066 13744 15092
rect 10176 14998 10202 15024
rect 12016 14998 12042 15024
rect 13396 14998 13422 15024
rect 14500 15121 14526 15126
rect 14500 15104 14515 15121
rect 14515 15104 14526 15121
rect 14822 15134 14848 15160
rect 15282 15134 15308 15160
rect 15604 15155 15630 15160
rect 15604 15138 15606 15155
rect 15606 15138 15630 15155
rect 15604 15134 15630 15138
rect 20756 15155 20782 15160
rect 20756 15138 20758 15155
rect 20758 15138 20782 15155
rect 20756 15134 20782 15138
rect 28392 15134 28418 15160
rect 28576 15134 28602 15160
rect 14500 15100 14526 15104
rect 15236 15100 15262 15126
rect 15512 15121 15538 15126
rect 15512 15104 15533 15121
rect 15533 15104 15538 15121
rect 15512 15100 15538 15104
rect 18410 15100 18436 15126
rect 18916 15121 18942 15126
rect 18916 15104 18920 15121
rect 18920 15104 18937 15121
rect 18937 15104 18942 15121
rect 18916 15100 18942 15104
rect 20250 15100 20276 15126
rect 20572 15100 20598 15126
rect 20802 15100 20828 15126
rect 28300 15100 28326 15126
rect 14270 15066 14296 15092
rect 15190 15066 15216 15092
rect 16018 14998 16044 15024
rect 28300 15032 28326 15058
rect 31750 15032 31776 15058
rect 29450 14998 29476 15024
rect 3322 14896 3348 14922
rect 3460 14896 3486 14922
rect 4840 14896 4866 14922
rect 6450 14896 6476 14922
rect 9210 14896 9236 14922
rect 10452 14862 10478 14888
rect 3184 14794 3210 14820
rect 5116 14828 5142 14854
rect 4794 14815 4820 14820
rect 4794 14798 4798 14815
rect 4798 14798 4815 14815
rect 4815 14798 4820 14815
rect 4794 14794 4820 14798
rect 4840 14794 4866 14820
rect 5898 14815 5924 14820
rect 5898 14798 5902 14815
rect 5902 14798 5919 14815
rect 5919 14798 5924 14815
rect 5898 14794 5924 14798
rect 6036 14815 6062 14820
rect 6036 14798 6057 14815
rect 6057 14798 6062 14815
rect 6036 14794 6062 14798
rect 3368 14781 3394 14786
rect 3368 14764 3370 14781
rect 3370 14764 3394 14781
rect 3368 14760 3394 14764
rect 4886 14781 4912 14786
rect 4886 14764 4890 14781
rect 4890 14764 4907 14781
rect 4907 14764 4912 14781
rect 4886 14760 4912 14764
rect 4932 14781 4958 14786
rect 4932 14764 4936 14781
rect 4936 14764 4953 14781
rect 4953 14764 4958 14781
rect 4932 14760 4958 14764
rect 6128 14781 6154 14786
rect 6128 14764 6130 14781
rect 6130 14764 6154 14781
rect 7002 14794 7028 14820
rect 7416 14815 7442 14820
rect 7416 14798 7420 14815
rect 7420 14798 7437 14815
rect 7437 14798 7442 14815
rect 7416 14794 7442 14798
rect 7462 14815 7488 14820
rect 7462 14798 7466 14815
rect 7466 14798 7483 14815
rect 7483 14798 7488 14815
rect 7462 14794 7488 14798
rect 7692 14794 7718 14820
rect 8290 14794 8316 14820
rect 6128 14760 6154 14764
rect 8244 14760 8270 14786
rect 8520 14794 8546 14820
rect 8934 14794 8960 14820
rect 8980 14794 9006 14820
rect 10176 14815 10202 14820
rect 10176 14798 10180 14815
rect 10180 14798 10197 14815
rect 10197 14798 10202 14815
rect 10176 14794 10202 14798
rect 8704 14760 8730 14786
rect 8888 14760 8914 14786
rect 12062 14896 12088 14922
rect 12568 14896 12594 14922
rect 13028 14896 13054 14922
rect 15788 14896 15814 14922
rect 16570 14896 16596 14922
rect 12292 14862 12318 14888
rect 10774 14828 10800 14854
rect 11418 14849 11444 14854
rect 11418 14832 11422 14849
rect 11422 14832 11439 14849
rect 11439 14832 11444 14849
rect 11418 14828 11444 14832
rect 13672 14862 13698 14888
rect 11694 14794 11720 14820
rect 11740 14794 11766 14820
rect 12292 14794 12318 14820
rect 13396 14815 13422 14820
rect 13396 14798 13400 14815
rect 13400 14798 13417 14815
rect 13417 14798 13422 14815
rect 13396 14794 13422 14798
rect 10544 14760 10570 14786
rect 13534 14813 13560 14820
rect 13534 14796 13551 14813
rect 13551 14796 13560 14813
rect 13810 14828 13836 14854
rect 14178 14849 14204 14854
rect 14178 14832 14182 14849
rect 14182 14832 14199 14849
rect 14199 14832 14204 14849
rect 14178 14828 14204 14832
rect 16018 14828 16044 14854
rect 24160 14828 24186 14854
rect 24344 14828 24370 14854
rect 13534 14794 13560 14796
rect 13718 14815 13744 14820
rect 13718 14798 13729 14815
rect 13729 14798 13744 14815
rect 13718 14794 13744 14798
rect 15880 14794 15906 14820
rect 21538 14794 21564 14820
rect 22044 14794 22070 14820
rect 24390 14794 24416 14820
rect 24758 14815 24784 14820
rect 24758 14798 24779 14815
rect 24779 14798 24784 14815
rect 24758 14794 24784 14798
rect 13810 14760 13836 14786
rect 13948 14760 13974 14786
rect 14224 14760 14250 14786
rect 14408 14781 14434 14786
rect 14408 14764 14410 14781
rect 14410 14764 14434 14781
rect 14408 14760 14434 14764
rect 16156 14760 16182 14786
rect 3184 14726 3210 14752
rect 5944 14726 5970 14752
rect 10176 14747 10202 14752
rect 10176 14730 10180 14747
rect 10180 14730 10197 14747
rect 10197 14730 10202 14747
rect 10176 14726 10202 14730
rect 10360 14726 10386 14752
rect 13902 14726 13928 14752
rect 16064 14747 16090 14752
rect 16064 14730 16068 14747
rect 16068 14730 16085 14747
rect 16085 14730 16090 14747
rect 16064 14726 16090 14730
rect 25908 14726 25934 14752
rect 4932 14624 4958 14650
rect 7462 14624 7488 14650
rect 11694 14624 11720 14650
rect 3828 14590 3854 14616
rect 9348 14611 9374 14616
rect 3184 14556 3210 14582
rect 3414 14556 3440 14582
rect 5898 14556 5924 14582
rect 3322 14522 3348 14548
rect 6818 14577 6844 14582
rect 6818 14560 6839 14577
rect 6839 14560 6844 14577
rect 9348 14594 9350 14611
rect 9350 14594 9374 14611
rect 9348 14590 9374 14594
rect 10268 14590 10294 14616
rect 11740 14590 11766 14616
rect 13534 14624 13560 14650
rect 12660 14590 12686 14616
rect 15420 14611 15446 14616
rect 15420 14594 15422 14611
rect 15422 14594 15446 14611
rect 15420 14590 15446 14594
rect 26460 14590 26486 14616
rect 6818 14556 6844 14560
rect 7094 14556 7120 14582
rect 8934 14556 8960 14582
rect 9256 14577 9282 14582
rect 9256 14560 9277 14577
rect 9277 14560 9282 14577
rect 9256 14556 9282 14560
rect 11418 14556 11444 14582
rect 12384 14577 12410 14582
rect 12384 14560 12388 14577
rect 12388 14560 12405 14577
rect 12405 14560 12410 14577
rect 12384 14556 12410 14560
rect 12522 14577 12548 14582
rect 12522 14560 12543 14577
rect 12543 14560 12548 14577
rect 12522 14556 12548 14560
rect 14224 14556 14250 14582
rect 15466 14556 15492 14582
rect 26138 14556 26164 14582
rect 28300 14556 28326 14582
rect 29358 14577 29384 14582
rect 29358 14560 29362 14577
rect 29362 14560 29379 14577
rect 29379 14560 29384 14577
rect 29358 14556 29384 14560
rect 29450 14577 29476 14582
rect 29450 14560 29454 14577
rect 29454 14560 29471 14577
rect 29471 14560 29476 14577
rect 29450 14556 29476 14560
rect 8520 14522 8546 14548
rect 9118 14543 9144 14548
rect 9118 14526 9122 14543
rect 9122 14526 9139 14543
rect 9139 14526 9144 14543
rect 9118 14522 9144 14526
rect 14178 14522 14204 14548
rect 15190 14543 15216 14548
rect 15190 14526 15194 14543
rect 15194 14526 15211 14543
rect 15211 14526 15216 14543
rect 15190 14522 15216 14526
rect 26000 14522 26026 14548
rect 6864 14454 6890 14480
rect 7278 14454 7304 14480
rect 10360 14454 10386 14480
rect 16202 14454 16228 14480
rect 22918 14454 22944 14480
rect 24298 14454 24324 14480
rect 27518 14454 27544 14480
rect 29588 14454 29614 14480
rect 3322 14352 3348 14378
rect 4978 14352 5004 14378
rect 6910 14352 6936 14378
rect 8842 14352 8868 14378
rect 4978 14284 5004 14310
rect 5254 14284 5280 14310
rect 5714 14284 5740 14310
rect 7278 14284 7304 14310
rect 7646 14305 7672 14310
rect 7646 14288 7650 14305
rect 7650 14288 7667 14305
rect 7667 14288 7672 14305
rect 7646 14284 7672 14288
rect 3184 14250 3210 14276
rect 3460 14250 3486 14276
rect 4794 14250 4820 14276
rect 5116 14250 5142 14276
rect 6036 14250 6062 14276
rect 6956 14250 6982 14276
rect 7784 14271 7810 14276
rect 7784 14254 7805 14271
rect 7805 14254 7810 14271
rect 7784 14250 7810 14254
rect 8704 14250 8730 14276
rect 10774 14250 10800 14276
rect 11004 14250 11030 14276
rect 11142 14250 11168 14276
rect 12154 14271 12180 14276
rect 12154 14254 12158 14271
rect 12158 14254 12175 14271
rect 12175 14254 12180 14271
rect 12154 14250 12180 14254
rect 12200 14271 12226 14276
rect 12200 14254 12204 14271
rect 12204 14254 12221 14271
rect 12221 14254 12226 14271
rect 12200 14250 12226 14254
rect 12384 14271 12410 14276
rect 12384 14254 12388 14271
rect 12388 14254 12405 14271
rect 12405 14254 12410 14271
rect 14500 14352 14526 14378
rect 15144 14352 15170 14378
rect 17168 14352 17194 14378
rect 22688 14352 22714 14378
rect 15650 14318 15676 14344
rect 21492 14318 21518 14344
rect 25816 14318 25842 14344
rect 25908 14318 25934 14344
rect 12384 14250 12410 14254
rect 13258 14271 13284 14276
rect 13258 14254 13262 14271
rect 13262 14254 13279 14271
rect 13279 14254 13284 14271
rect 13258 14250 13284 14254
rect 11096 14237 11122 14242
rect 11096 14220 11098 14237
rect 11098 14220 11122 14237
rect 11096 14216 11122 14220
rect 12292 14237 12318 14242
rect 12292 14220 12296 14237
rect 12296 14220 12313 14237
rect 12313 14220 12318 14237
rect 12292 14216 12318 14220
rect 12246 14203 12272 14208
rect 12246 14186 12250 14203
rect 12250 14186 12267 14203
rect 12267 14186 12272 14203
rect 12246 14182 12272 14186
rect 12338 14182 12364 14208
rect 13810 14250 13836 14276
rect 17674 14271 17700 14276
rect 17674 14254 17678 14271
rect 17678 14254 17695 14271
rect 17695 14254 17700 14271
rect 17674 14250 17700 14254
rect 17904 14284 17930 14310
rect 19284 14284 19310 14310
rect 21354 14305 21380 14310
rect 21354 14288 21358 14305
rect 21358 14288 21375 14305
rect 21375 14288 21380 14305
rect 21354 14284 21380 14288
rect 24344 14305 24370 14310
rect 24344 14288 24348 14305
rect 24348 14288 24365 14305
rect 24365 14288 24370 14305
rect 24344 14284 24370 14288
rect 19376 14250 19402 14276
rect 19882 14250 19908 14276
rect 21124 14250 21150 14276
rect 22872 14271 22898 14276
rect 22872 14254 22876 14271
rect 22876 14254 22893 14271
rect 22893 14254 22898 14271
rect 22872 14250 22898 14254
rect 24666 14250 24692 14276
rect 25632 14271 25658 14276
rect 25632 14254 25636 14271
rect 25636 14254 25653 14271
rect 25653 14254 25658 14271
rect 25632 14250 25658 14254
rect 25770 14271 25796 14276
rect 25770 14254 25787 14271
rect 25787 14254 25796 14271
rect 25770 14250 25796 14254
rect 28254 14352 28280 14378
rect 26000 14250 26026 14276
rect 27702 14271 27728 14276
rect 27702 14254 27706 14271
rect 27706 14254 27723 14271
rect 27723 14254 27728 14271
rect 27702 14250 27728 14254
rect 17766 14216 17792 14242
rect 23102 14216 23128 14242
rect 24390 14216 24416 14242
rect 24574 14237 24600 14242
rect 24574 14220 24576 14237
rect 24576 14220 24600 14237
rect 24574 14216 24600 14220
rect 28346 14250 28372 14276
rect 28438 14250 28464 14276
rect 17214 14182 17240 14208
rect 17720 14203 17746 14208
rect 17720 14186 17724 14203
rect 17724 14186 17741 14203
rect 17741 14186 17746 14203
rect 17720 14182 17746 14186
rect 17812 14203 17838 14208
rect 17812 14186 17816 14203
rect 17816 14186 17833 14203
rect 17833 14186 17838 14203
rect 17812 14182 17838 14186
rect 19514 14203 19540 14208
rect 19514 14186 19518 14203
rect 19518 14186 19535 14203
rect 19535 14186 19540 14203
rect 19514 14182 19540 14186
rect 21446 14182 21472 14208
rect 26828 14182 26854 14208
rect 28576 14182 28602 14208
rect 11096 14080 11122 14106
rect 14454 14080 14480 14106
rect 17766 14101 17792 14106
rect 17766 14084 17770 14101
rect 17770 14084 17787 14101
rect 17787 14084 17792 14101
rect 17766 14080 17792 14084
rect 19882 14080 19908 14106
rect 3184 14046 3210 14072
rect 4794 14012 4820 14038
rect 5254 14012 5280 14038
rect 6404 14046 6430 14072
rect 12292 14046 12318 14072
rect 3322 13978 3348 14004
rect 6266 14033 6292 14038
rect 6266 14016 6270 14033
rect 6270 14016 6287 14033
rect 6287 14016 6292 14033
rect 6266 14012 6292 14016
rect 6450 14012 6476 14038
rect 9624 14033 9650 14038
rect 9624 14016 9628 14033
rect 9628 14016 9645 14033
rect 9645 14016 9650 14033
rect 9624 14012 9650 14016
rect 9762 14033 9788 14038
rect 9762 14016 9766 14033
rect 9766 14016 9783 14033
rect 9783 14016 9788 14033
rect 9762 14012 9788 14016
rect 6312 13944 6338 13970
rect 17260 14046 17286 14072
rect 19376 14046 19402 14072
rect 20618 14080 20644 14106
rect 21354 14080 21380 14106
rect 21446 14101 21472 14106
rect 21446 14084 21450 14101
rect 21450 14084 21467 14101
rect 21467 14084 21472 14101
rect 21446 14080 21472 14084
rect 22826 14080 22852 14106
rect 24114 14080 24140 14106
rect 25816 14080 25842 14106
rect 15328 14012 15354 14038
rect 15190 13978 15216 14004
rect 15420 14033 15446 14038
rect 15420 14016 15424 14033
rect 15424 14016 15441 14033
rect 15441 14016 15446 14033
rect 15420 14012 15446 14016
rect 15650 14012 15676 14038
rect 16754 14012 16780 14038
rect 17674 14012 17700 14038
rect 19882 14033 19908 14038
rect 19882 14016 19886 14033
rect 19886 14016 19903 14033
rect 19903 14016 19908 14033
rect 19882 14012 19908 14016
rect 19974 14012 20000 14038
rect 21492 14046 21518 14072
rect 26184 14067 26210 14072
rect 26184 14050 26186 14067
rect 26186 14050 26210 14067
rect 26184 14046 26210 14050
rect 16938 13978 16964 14004
rect 17076 13999 17102 14004
rect 17076 13982 17080 13999
rect 17080 13982 17097 13999
rect 17097 13982 17102 13999
rect 17076 13978 17102 13982
rect 20066 13999 20092 14004
rect 20066 13982 20070 13999
rect 20070 13982 20087 13999
rect 20087 13982 20092 13999
rect 20066 13978 20092 13982
rect 20802 13978 20828 14004
rect 12384 13944 12410 13970
rect 21492 13978 21518 14004
rect 5208 13910 5234 13936
rect 6404 13931 6430 13936
rect 6404 13914 6408 13931
rect 6408 13914 6425 13931
rect 6425 13914 6430 13931
rect 6404 13910 6430 13914
rect 9670 13910 9696 13936
rect 14592 13910 14618 13936
rect 20066 13910 20092 13936
rect 20618 13910 20644 13936
rect 22918 13910 22944 13936
rect 24390 14012 24416 14038
rect 26092 14033 26118 14038
rect 27426 14080 27452 14106
rect 27518 14080 27544 14106
rect 26092 14016 26113 14033
rect 26113 14016 26118 14033
rect 26092 14012 26118 14016
rect 25954 13999 25980 14004
rect 25954 13982 25958 13999
rect 25958 13982 25975 13999
rect 25975 13982 25980 13999
rect 25954 13978 25980 13982
rect 27104 13978 27130 14004
rect 27393 14033 27419 14038
rect 27393 14016 27397 14033
rect 27397 14016 27414 14033
rect 27414 14016 27419 14033
rect 27393 14012 27419 14016
rect 27564 14033 27590 14038
rect 27564 14016 27575 14033
rect 27575 14016 27590 14033
rect 27564 14012 27590 14016
rect 28254 14033 28280 14038
rect 28254 14016 28275 14033
rect 28275 14016 28280 14033
rect 28254 14012 28280 14016
rect 28438 14012 28464 14038
rect 27150 13944 27176 13970
rect 27288 13944 27314 13970
rect 27702 13978 27728 14004
rect 28070 13978 28096 14004
rect 26230 13910 26256 13936
rect 27242 13931 27268 13936
rect 27242 13914 27246 13931
rect 27246 13914 27263 13931
rect 27263 13914 27268 13931
rect 27242 13910 27268 13914
rect 28990 13910 29016 13936
rect 6266 13808 6292 13834
rect 9624 13808 9650 13834
rect 7646 13740 7672 13766
rect 8474 13761 8500 13766
rect 8474 13744 8478 13761
rect 8478 13744 8495 13761
rect 8495 13744 8500 13761
rect 8474 13740 8500 13744
rect 5208 13706 5234 13732
rect 5714 13706 5740 13732
rect 8612 13706 8638 13732
rect 8888 13706 8914 13732
rect 10038 13706 10064 13732
rect 10774 13808 10800 13834
rect 12200 13808 12226 13834
rect 15420 13808 15446 13834
rect 16754 13829 16780 13834
rect 16754 13812 16758 13829
rect 16758 13812 16775 13829
rect 16775 13812 16780 13829
rect 16754 13808 16780 13812
rect 22320 13808 22346 13834
rect 22688 13808 22714 13834
rect 25770 13808 25796 13834
rect 27058 13808 27084 13834
rect 27564 13808 27590 13834
rect 24068 13774 24094 13800
rect 25356 13774 25382 13800
rect 16800 13761 16826 13766
rect 16800 13744 16804 13761
rect 16804 13744 16821 13761
rect 16821 13744 16826 13761
rect 16800 13740 16826 13744
rect 17076 13740 17102 13766
rect 24344 13740 24370 13766
rect 10728 13706 10754 13732
rect 11004 13706 11030 13732
rect 14178 13727 14204 13732
rect 14178 13710 14182 13727
rect 14182 13710 14199 13727
rect 14199 13710 14204 13727
rect 14178 13706 14204 13710
rect 5116 13672 5142 13698
rect 5392 13693 5418 13698
rect 5392 13676 5394 13693
rect 5394 13676 5418 13693
rect 5392 13672 5418 13676
rect 8750 13672 8776 13698
rect 10912 13693 10938 13698
rect 10912 13676 10914 13693
rect 10914 13676 10938 13693
rect 10912 13672 10938 13676
rect 12936 13672 12962 13698
rect 14500 13706 14526 13732
rect 15926 13706 15952 13732
rect 17812 13706 17838 13732
rect 23102 13727 23128 13732
rect 23102 13710 23106 13727
rect 23106 13710 23123 13727
rect 23123 13710 23128 13727
rect 23102 13706 23128 13710
rect 23148 13727 23174 13732
rect 23148 13710 23152 13727
rect 23152 13710 23169 13727
rect 23169 13710 23174 13727
rect 23148 13706 23174 13710
rect 24390 13706 24416 13732
rect 26828 13727 26854 13732
rect 26828 13710 26832 13727
rect 26832 13710 26849 13727
rect 26849 13710 26854 13727
rect 26828 13706 26854 13710
rect 27242 13740 27268 13766
rect 27150 13706 27176 13732
rect 14454 13672 14480 13698
rect 18824 13693 18850 13698
rect 18824 13676 18841 13693
rect 18841 13676 18850 13693
rect 18824 13672 18850 13676
rect 21492 13672 21518 13698
rect 24712 13693 24738 13698
rect 24712 13676 24714 13693
rect 24714 13676 24738 13693
rect 24712 13672 24738 13676
rect 28898 13706 28924 13732
rect 29496 13727 29522 13732
rect 29496 13710 29500 13727
rect 29500 13710 29517 13727
rect 29517 13710 29522 13727
rect 29496 13706 29522 13710
rect 29588 13727 29614 13732
rect 29588 13710 29592 13727
rect 29592 13710 29609 13727
rect 29609 13710 29614 13727
rect 29588 13706 29614 13710
rect 19376 13659 19402 13664
rect 19376 13642 19380 13659
rect 19380 13642 19397 13659
rect 19397 13642 19402 13659
rect 19376 13638 19402 13642
rect 28576 13672 28602 13698
rect 28714 13693 28740 13698
rect 28714 13676 28718 13693
rect 28718 13676 28735 13693
rect 28735 13676 28740 13693
rect 28714 13672 28740 13676
rect 28990 13672 29016 13698
rect 29542 13659 29568 13664
rect 29542 13642 29546 13659
rect 29546 13642 29563 13659
rect 29563 13642 29568 13659
rect 29542 13638 29568 13642
rect 5024 13536 5050 13562
rect 9670 13557 9696 13562
rect 9670 13540 9674 13557
rect 9674 13540 9691 13557
rect 9691 13540 9696 13557
rect 9670 13536 9696 13540
rect 15328 13536 15354 13562
rect 16294 13557 16320 13562
rect 16294 13540 16298 13557
rect 16298 13540 16315 13557
rect 16315 13540 16320 13557
rect 16294 13536 16320 13540
rect 3552 13523 3578 13528
rect 3552 13506 3554 13523
rect 3554 13506 3578 13523
rect 3552 13502 3578 13506
rect 6956 13502 6982 13528
rect 7186 13502 7212 13528
rect 8290 13502 8316 13528
rect 9854 13502 9880 13528
rect 10268 13523 10294 13528
rect 10268 13506 10270 13523
rect 10270 13506 10294 13523
rect 10268 13502 10294 13506
rect 11648 13502 11674 13528
rect 14546 13523 14572 13528
rect 14546 13506 14548 13523
rect 14548 13506 14572 13523
rect 3322 13489 3348 13494
rect 3322 13472 3326 13489
rect 3326 13472 3343 13489
rect 3343 13472 3348 13489
rect 3322 13468 3348 13472
rect 3460 13489 3486 13494
rect 3460 13472 3481 13489
rect 3481 13472 3486 13489
rect 3460 13468 3486 13472
rect 4610 13489 4636 13494
rect 4610 13472 4614 13489
rect 4614 13472 4631 13489
rect 4631 13472 4636 13489
rect 4610 13468 4636 13472
rect 5024 13468 5050 13494
rect 5162 13489 5188 13494
rect 5162 13472 5166 13489
rect 5166 13472 5183 13489
rect 5183 13472 5188 13489
rect 5162 13468 5188 13472
rect 6312 13468 6338 13494
rect 6864 13434 6890 13460
rect 9256 13489 9282 13494
rect 9256 13472 9260 13489
rect 9260 13472 9277 13489
rect 9277 13472 9282 13489
rect 9256 13468 9282 13472
rect 10314 13468 10340 13494
rect 10728 13468 10754 13494
rect 5116 13400 5142 13426
rect 6174 13366 6200 13392
rect 8106 13400 8132 13426
rect 10038 13455 10064 13460
rect 10038 13438 10042 13455
rect 10042 13438 10059 13455
rect 10059 13438 10064 13455
rect 10038 13434 10064 13438
rect 8014 13366 8040 13392
rect 9946 13366 9972 13392
rect 12430 13489 12456 13494
rect 12430 13472 12434 13489
rect 12434 13472 12451 13489
rect 12451 13472 12456 13489
rect 12430 13468 12456 13472
rect 12522 13468 12548 13494
rect 12936 13489 12962 13494
rect 12936 13472 12957 13489
rect 12957 13472 12962 13489
rect 14546 13502 14572 13506
rect 12936 13468 12962 13472
rect 14362 13468 14388 13494
rect 14454 13489 14480 13494
rect 14454 13472 14475 13489
rect 14475 13472 14480 13489
rect 14454 13468 14480 13472
rect 17076 13502 17102 13528
rect 17720 13502 17746 13528
rect 17858 13502 17884 13528
rect 19376 13536 19402 13562
rect 27426 13536 27452 13562
rect 16018 13468 16044 13494
rect 18318 13468 18344 13494
rect 19514 13502 19540 13528
rect 19054 13489 19080 13494
rect 19054 13472 19058 13489
rect 19058 13472 19075 13489
rect 19075 13472 19080 13489
rect 19054 13468 19080 13472
rect 25356 13468 25382 13494
rect 26000 13489 26026 13494
rect 26000 13472 26004 13489
rect 26004 13472 26021 13489
rect 26021 13472 26026 13489
rect 26000 13468 26026 13472
rect 26138 13489 26164 13494
rect 26138 13472 26159 13489
rect 26159 13472 26164 13489
rect 26138 13468 26164 13472
rect 26322 13468 26348 13494
rect 27012 13468 27038 13494
rect 12752 13434 12778 13460
rect 12798 13455 12824 13460
rect 12798 13438 12802 13455
rect 12802 13438 12819 13455
rect 12819 13438 12824 13455
rect 12798 13434 12824 13438
rect 14178 13434 14204 13460
rect 14316 13455 14342 13460
rect 14316 13438 14320 13455
rect 14320 13438 14337 13455
rect 14337 13438 14342 13455
rect 14316 13434 14342 13438
rect 15604 13455 15630 13460
rect 15604 13438 15608 13455
rect 15608 13438 15625 13455
rect 15625 13438 15630 13455
rect 15604 13434 15630 13438
rect 20066 13434 20092 13460
rect 21400 13434 21426 13460
rect 21584 13434 21610 13460
rect 24160 13455 24186 13460
rect 24160 13438 24164 13455
rect 24164 13438 24181 13455
rect 24181 13438 24186 13455
rect 24160 13434 24186 13438
rect 18732 13400 18758 13426
rect 18778 13400 18804 13426
rect 21354 13400 21380 13426
rect 11878 13366 11904 13392
rect 12476 13366 12502 13392
rect 14684 13366 14710 13392
rect 16524 13366 16550 13392
rect 24252 13387 24278 13392
rect 24252 13370 24256 13387
rect 24256 13370 24273 13387
rect 24273 13370 24278 13387
rect 24252 13366 24278 13370
rect 3322 13264 3348 13290
rect 4610 13264 4636 13290
rect 4840 13264 4866 13290
rect 8198 13264 8224 13290
rect 10084 13264 10110 13290
rect 8290 13230 8316 13256
rect 3138 13217 3164 13222
rect 3138 13200 3142 13217
rect 3142 13200 3159 13217
rect 3159 13200 3164 13217
rect 3138 13196 3164 13200
rect 5162 13196 5188 13222
rect 5208 13196 5234 13222
rect 5346 13217 5372 13222
rect 5346 13200 5350 13217
rect 5350 13200 5367 13217
rect 5367 13200 5372 13217
rect 5346 13196 5372 13200
rect 3460 13162 3486 13188
rect 4748 13183 4774 13188
rect 4748 13166 4752 13183
rect 4752 13166 4769 13183
rect 4769 13166 4774 13183
rect 4748 13162 4774 13166
rect 4840 13183 4866 13188
rect 4840 13166 4847 13183
rect 4847 13166 4864 13183
rect 4864 13166 4866 13183
rect 4840 13162 4866 13166
rect 5392 13162 5418 13188
rect 3368 13149 3394 13154
rect 3368 13132 3370 13149
rect 3370 13132 3394 13149
rect 3368 13128 3394 13132
rect 4656 13149 4682 13154
rect 4656 13132 4660 13149
rect 4660 13132 4677 13149
rect 4677 13132 4682 13149
rect 4656 13128 4682 13132
rect 4794 13149 4820 13154
rect 4794 13132 4798 13149
rect 4798 13132 4815 13149
rect 4815 13132 4820 13149
rect 4794 13128 4820 13132
rect 5300 13128 5326 13154
rect 7876 13183 7902 13188
rect 7876 13166 7880 13183
rect 7880 13166 7897 13183
rect 7897 13166 7902 13183
rect 7876 13162 7902 13166
rect 7922 13183 7948 13188
rect 7922 13166 7937 13183
rect 7937 13166 7948 13183
rect 7922 13162 7948 13166
rect 8014 13181 8040 13188
rect 8014 13164 8031 13181
rect 8031 13164 8040 13181
rect 8014 13162 8040 13164
rect 8089 13183 8115 13188
rect 8089 13166 8093 13183
rect 8093 13166 8110 13183
rect 8110 13166 8115 13183
rect 8089 13162 8115 13166
rect 8198 13183 8224 13188
rect 8198 13166 8209 13183
rect 8209 13166 8224 13183
rect 8198 13162 8224 13166
rect 8474 13162 8500 13188
rect 10038 13196 10064 13222
rect 12430 13264 12456 13290
rect 12752 13264 12778 13290
rect 14684 13230 14710 13256
rect 8612 13128 8638 13154
rect 11050 13162 11076 13188
rect 11004 13128 11030 13154
rect 12798 13162 12824 13188
rect 13580 13162 13606 13188
rect 14500 13162 14526 13188
rect 14638 13183 14664 13188
rect 14638 13166 14644 13183
rect 14644 13166 14664 13183
rect 14638 13162 14664 13166
rect 15880 13264 15906 13290
rect 16018 13264 16044 13290
rect 18824 13264 18850 13290
rect 24160 13264 24186 13290
rect 29542 13264 29568 13290
rect 14822 13230 14848 13256
rect 23148 13230 23174 13256
rect 28760 13230 28786 13256
rect 16938 13196 16964 13222
rect 11280 13128 11306 13154
rect 11648 13149 11674 13154
rect 11648 13132 11650 13149
rect 11650 13132 11674 13149
rect 11648 13128 11674 13132
rect 12936 13128 12962 13154
rect 14960 13162 14986 13188
rect 16294 13162 16320 13188
rect 16570 13162 16596 13188
rect 18686 13162 18712 13188
rect 18732 13183 18758 13188
rect 18732 13166 18736 13183
rect 18736 13166 18753 13183
rect 18753 13166 18758 13183
rect 18732 13162 18758 13166
rect 20848 13196 20874 13222
rect 21216 13183 21242 13188
rect 21216 13166 21220 13183
rect 21220 13166 21237 13183
rect 21237 13166 21242 13183
rect 21216 13162 21242 13166
rect 21538 13162 21564 13188
rect 21906 13162 21932 13188
rect 22826 13162 22852 13188
rect 6358 13094 6384 13120
rect 8152 13094 8178 13120
rect 9762 13094 9788 13120
rect 14546 13115 14572 13120
rect 14546 13098 14550 13115
rect 14550 13098 14567 13115
rect 14567 13098 14572 13115
rect 14546 13094 14572 13098
rect 19284 13128 19310 13154
rect 14822 13094 14848 13120
rect 17168 13094 17194 13120
rect 22872 13094 22898 13120
rect 4794 12992 4820 13018
rect 5300 12992 5326 13018
rect 5622 12992 5648 13018
rect 8152 12992 8178 13018
rect 12384 13013 12410 13018
rect 12384 12996 12388 13013
rect 12388 12996 12405 13013
rect 12405 12996 12410 13013
rect 12384 12992 12410 12996
rect 14500 12992 14526 13018
rect 19284 12992 19310 13018
rect 22780 12992 22806 13018
rect 3874 12979 3900 12984
rect 3874 12962 3876 12979
rect 3876 12962 3900 12979
rect 3874 12958 3900 12962
rect 3460 12924 3486 12950
rect 3920 12924 3946 12950
rect 6312 12979 6338 12984
rect 6312 12962 6316 12979
rect 6316 12962 6333 12979
rect 6333 12962 6338 12979
rect 6312 12958 6338 12962
rect 6358 12979 6384 12984
rect 6358 12962 6362 12979
rect 6362 12962 6379 12979
rect 6379 12962 6384 12979
rect 6358 12958 6384 12962
rect 3138 12890 3164 12916
rect 6174 12945 6200 12950
rect 6174 12928 6178 12945
rect 6178 12928 6195 12945
rect 6195 12928 6200 12945
rect 6174 12924 6200 12928
rect 6220 12945 6246 12950
rect 6220 12928 6224 12945
rect 6224 12928 6241 12945
rect 6241 12928 6246 12945
rect 6220 12924 6246 12928
rect 6450 12958 6476 12984
rect 6496 12890 6522 12916
rect 7094 12945 7120 12950
rect 7094 12928 7115 12945
rect 7115 12928 7120 12945
rect 10084 12958 10110 12984
rect 13028 12979 13054 12984
rect 7094 12924 7120 12928
rect 9118 12924 9144 12950
rect 10314 12924 10340 12950
rect 11740 12945 11766 12950
rect 11740 12928 11744 12945
rect 11744 12928 11761 12945
rect 11761 12928 11766 12945
rect 11740 12924 11766 12928
rect 13028 12962 13030 12979
rect 13030 12962 13054 12979
rect 13028 12958 13054 12962
rect 11878 12945 11904 12950
rect 11878 12928 11895 12945
rect 11895 12928 11904 12945
rect 12062 12945 12088 12950
rect 11878 12924 11904 12928
rect 12062 12928 12073 12945
rect 12073 12928 12088 12945
rect 12062 12924 12088 12928
rect 12246 12924 12272 12950
rect 12476 12945 12502 12950
rect 12476 12928 12480 12945
rect 12480 12928 12497 12945
rect 12497 12928 12502 12945
rect 12476 12924 12502 12928
rect 12936 12945 12962 12950
rect 16432 12958 16458 12984
rect 17444 12958 17470 12984
rect 19238 12979 19264 12984
rect 19238 12962 19242 12979
rect 19242 12962 19259 12979
rect 19259 12962 19264 12979
rect 19238 12958 19264 12962
rect 12936 12928 12957 12945
rect 12957 12928 12962 12945
rect 12936 12924 12962 12928
rect 16478 12945 16504 12950
rect 16478 12928 16482 12945
rect 16482 12928 16499 12945
rect 16499 12928 16504 12945
rect 16478 12924 16504 12928
rect 20802 12958 20828 12984
rect 20848 12958 20874 12984
rect 21032 12979 21058 12984
rect 21032 12962 21034 12979
rect 21034 12962 21058 12979
rect 21032 12958 21058 12962
rect 22826 12958 22852 12984
rect 19376 12945 19402 12950
rect 19376 12928 19380 12945
rect 19380 12928 19397 12945
rect 19397 12928 19402 12945
rect 19376 12924 19402 12928
rect 22642 12945 22668 12950
rect 22642 12928 22657 12945
rect 22657 12928 22668 12945
rect 22642 12924 22668 12928
rect 6864 12822 6890 12848
rect 10038 12911 10064 12916
rect 10038 12894 10042 12911
rect 10042 12894 10059 12911
rect 10059 12894 10064 12911
rect 10038 12890 10064 12894
rect 9026 12822 9052 12848
rect 10268 12822 10294 12848
rect 12798 12911 12824 12916
rect 12798 12894 12802 12911
rect 12802 12894 12819 12911
rect 12819 12894 12824 12911
rect 12798 12890 12824 12894
rect 16570 12890 16596 12916
rect 17076 12890 17102 12916
rect 19284 12911 19310 12916
rect 19284 12894 19288 12911
rect 19288 12894 19305 12911
rect 19305 12894 19310 12911
rect 19284 12890 19310 12894
rect 12062 12856 12088 12882
rect 12430 12843 12456 12848
rect 12430 12826 12434 12843
rect 12434 12826 12451 12843
rect 12451 12826 12456 12843
rect 12430 12822 12456 12826
rect 14822 12822 14848 12848
rect 22274 12890 22300 12916
rect 29496 13013 29522 13018
rect 29496 12996 29500 13013
rect 29500 12996 29517 13013
rect 29517 12996 29522 13013
rect 29496 12992 29522 12996
rect 25862 12958 25888 12984
rect 28116 12958 28142 12984
rect 28254 12958 28280 12984
rect 22918 12945 22944 12950
rect 22918 12928 22929 12945
rect 22929 12928 22944 12945
rect 22918 12924 22944 12928
rect 25632 12924 25658 12950
rect 26138 12924 26164 12950
rect 28530 12924 28556 12950
rect 29404 12924 29430 12950
rect 29542 12945 29568 12950
rect 29542 12928 29557 12945
rect 29557 12928 29568 12945
rect 29542 12924 29568 12928
rect 29634 12924 29660 12950
rect 29709 12945 29735 12950
rect 29709 12928 29713 12945
rect 29713 12928 29730 12945
rect 29730 12928 29735 12945
rect 29709 12924 29735 12928
rect 29818 12945 29844 12950
rect 29818 12928 29829 12945
rect 29829 12928 29844 12945
rect 22872 12856 22898 12882
rect 21216 12822 21242 12848
rect 22596 12843 22622 12848
rect 22596 12826 22600 12843
rect 22600 12826 22617 12843
rect 22617 12826 22622 12843
rect 22596 12822 22622 12826
rect 25540 12822 25566 12848
rect 27840 12890 27866 12916
rect 28070 12890 28096 12916
rect 29818 12924 29844 12928
rect 26000 12822 26026 12848
rect 27334 12822 27360 12848
rect 4656 12720 4682 12746
rect 3138 12673 3164 12678
rect 3138 12656 3142 12673
rect 3142 12656 3159 12673
rect 3159 12656 3164 12673
rect 3138 12652 3164 12656
rect 5346 12720 5372 12746
rect 6220 12720 6246 12746
rect 3460 12618 3486 12644
rect 5254 12618 5280 12644
rect 8336 12720 8362 12746
rect 9256 12720 9282 12746
rect 11280 12720 11306 12746
rect 12062 12720 12088 12746
rect 14040 12720 14066 12746
rect 22274 12720 22300 12746
rect 29542 12720 29568 12746
rect 6864 12652 6890 12678
rect 10038 12652 10064 12678
rect 6496 12639 6522 12644
rect 6496 12622 6500 12639
rect 6500 12622 6517 12639
rect 6517 12622 6522 12639
rect 6496 12618 6522 12622
rect 7232 12618 7258 12644
rect 10314 12618 10340 12644
rect 10452 12618 10478 12644
rect 3414 12584 3440 12610
rect 4748 12584 4774 12610
rect 4978 12584 5004 12610
rect 7416 12584 7442 12610
rect 8152 12584 8178 12610
rect 8336 12605 8362 12610
rect 8336 12588 8338 12605
rect 8338 12588 8362 12605
rect 8336 12584 8362 12588
rect 9118 12584 9144 12610
rect 13028 12618 13054 12644
rect 14592 12652 14618 12678
rect 14546 12639 14572 12644
rect 14546 12622 14550 12639
rect 14550 12622 14567 12639
rect 14567 12622 14572 12639
rect 14546 12618 14572 12622
rect 14684 12639 14710 12644
rect 14684 12622 14688 12639
rect 14688 12622 14705 12639
rect 14705 12622 14710 12639
rect 14684 12618 14710 12622
rect 15696 12639 15722 12644
rect 15696 12622 15700 12639
rect 15700 12622 15717 12639
rect 15717 12622 15722 12639
rect 15696 12618 15722 12622
rect 16570 12652 16596 12678
rect 19882 12652 19908 12678
rect 16432 12639 16458 12644
rect 16432 12622 16436 12639
rect 16436 12622 16453 12639
rect 16453 12622 16458 12639
rect 16432 12618 16458 12622
rect 16524 12639 16550 12644
rect 16524 12622 16528 12639
rect 16528 12622 16545 12639
rect 16545 12622 16550 12639
rect 16524 12618 16550 12622
rect 13902 12605 13928 12610
rect 13902 12588 13906 12605
rect 13906 12588 13923 12605
rect 13923 12588 13928 12605
rect 13902 12584 13928 12588
rect 16294 12584 16320 12610
rect 16478 12584 16504 12610
rect 19514 12618 19540 12644
rect 19974 12618 20000 12644
rect 21216 12673 21242 12678
rect 21216 12656 21220 12673
rect 21220 12656 21237 12673
rect 21237 12656 21242 12673
rect 21216 12652 21242 12656
rect 22412 12652 22438 12678
rect 22642 12652 22668 12678
rect 25586 12652 25612 12678
rect 26276 12652 26302 12678
rect 20434 12605 20460 12610
rect 20434 12588 20438 12605
rect 20438 12588 20455 12605
rect 20455 12588 20460 12605
rect 20434 12584 20460 12588
rect 20480 12584 20506 12610
rect 20848 12618 20874 12644
rect 21630 12618 21656 12644
rect 27840 12639 27866 12644
rect 27840 12622 27844 12639
rect 27844 12622 27861 12639
rect 27861 12622 27866 12639
rect 27840 12618 27866 12622
rect 28116 12618 28142 12644
rect 28162 12618 28188 12644
rect 28070 12605 28096 12610
rect 28070 12588 28072 12605
rect 28072 12588 28096 12605
rect 28070 12584 28096 12588
rect 3920 12550 3946 12576
rect 5254 12550 5280 12576
rect 6542 12571 6568 12576
rect 6542 12554 6546 12571
rect 6546 12554 6563 12571
rect 6563 12554 6568 12571
rect 6542 12550 6568 12554
rect 11694 12550 11720 12576
rect 12614 12550 12640 12576
rect 13994 12571 14020 12576
rect 13994 12554 14006 12571
rect 14006 12554 14020 12571
rect 13994 12550 14020 12554
rect 14730 12550 14756 12576
rect 15742 12571 15768 12576
rect 15742 12554 15746 12571
rect 15746 12554 15763 12571
rect 15763 12554 15768 12571
rect 15742 12550 15768 12554
rect 17168 12550 17194 12576
rect 18318 12550 18344 12576
rect 28300 12550 28326 12576
rect 28392 12550 28418 12576
rect 5254 12448 5280 12474
rect 5622 12448 5648 12474
rect 5944 12448 5970 12474
rect 10406 12448 10432 12474
rect 11694 12448 11720 12474
rect 3138 12414 3164 12440
rect 4748 12435 4774 12440
rect 4748 12418 4750 12435
rect 4750 12418 4774 12435
rect 4748 12414 4774 12418
rect 6910 12414 6936 12440
rect 8152 12414 8178 12440
rect 8612 12414 8638 12440
rect 9026 12435 9052 12440
rect 9026 12418 9028 12435
rect 9028 12418 9052 12435
rect 9026 12414 9052 12418
rect 12384 12448 12410 12474
rect 14822 12448 14848 12474
rect 16340 12448 16366 12474
rect 6542 12380 6568 12406
rect 6864 12401 6890 12406
rect 6864 12384 6868 12401
rect 6868 12384 6885 12401
rect 6885 12384 6890 12401
rect 6864 12380 6890 12384
rect 7140 12380 7166 12406
rect 7876 12380 7902 12406
rect 8474 12380 8500 12406
rect 10038 12380 10064 12406
rect 11556 12401 11582 12406
rect 11556 12384 11560 12401
rect 11560 12384 11577 12401
rect 11577 12384 11582 12401
rect 11556 12380 11582 12384
rect 4518 12367 4544 12372
rect 4518 12350 4522 12367
rect 4522 12350 4539 12367
rect 4539 12350 4544 12367
rect 4518 12346 4544 12350
rect 10866 12367 10892 12372
rect 10866 12350 10870 12367
rect 10870 12350 10887 12367
rect 10887 12350 10892 12367
rect 10866 12346 10892 12350
rect 12016 12435 12042 12440
rect 12016 12418 12020 12435
rect 12020 12418 12037 12435
rect 12037 12418 12042 12435
rect 12016 12414 12042 12418
rect 12614 12414 12640 12440
rect 11648 12401 11674 12406
rect 11648 12384 11652 12401
rect 11652 12384 11669 12401
rect 11669 12384 11674 12401
rect 11648 12380 11674 12384
rect 11694 12401 11720 12406
rect 11694 12384 11698 12401
rect 11698 12384 11715 12401
rect 11715 12384 11720 12401
rect 11694 12380 11720 12384
rect 11740 12401 11766 12406
rect 11740 12384 11747 12401
rect 11747 12384 11764 12401
rect 11764 12384 11766 12401
rect 11740 12380 11766 12384
rect 12890 12380 12916 12406
rect 14592 12414 14618 12440
rect 15742 12435 15768 12440
rect 15742 12418 15759 12435
rect 15759 12418 15768 12435
rect 15742 12414 15768 12418
rect 17076 12435 17102 12440
rect 17076 12418 17080 12435
rect 17080 12418 17097 12435
rect 17097 12418 17102 12435
rect 17076 12414 17102 12418
rect 15604 12401 15630 12406
rect 15604 12384 15608 12401
rect 15608 12384 15625 12401
rect 15625 12384 15630 12401
rect 15604 12380 15630 12384
rect 17030 12380 17056 12406
rect 17168 12401 17194 12406
rect 17168 12384 17172 12401
rect 17172 12384 17189 12401
rect 17189 12384 17194 12401
rect 17168 12380 17194 12384
rect 17214 12401 17240 12406
rect 17214 12384 17218 12401
rect 17218 12384 17235 12401
rect 17235 12384 17240 12401
rect 17214 12380 17240 12384
rect 5438 12278 5464 12304
rect 8934 12278 8960 12304
rect 11970 12278 11996 12304
rect 14316 12367 14342 12372
rect 14316 12350 14320 12367
rect 14320 12350 14337 12367
rect 14337 12350 14342 12367
rect 14316 12346 14342 12350
rect 12798 12278 12824 12304
rect 17214 12312 17240 12338
rect 17674 12380 17700 12406
rect 17858 12401 17884 12406
rect 17858 12384 17862 12401
rect 17862 12384 17879 12401
rect 17879 12384 17884 12401
rect 17858 12380 17884 12384
rect 17904 12401 17930 12406
rect 17904 12384 17908 12401
rect 17908 12384 17925 12401
rect 17925 12384 17930 12401
rect 17904 12380 17930 12384
rect 18318 12435 18344 12440
rect 18318 12418 18322 12435
rect 18322 12418 18339 12435
rect 18339 12418 18344 12435
rect 18318 12414 18344 12418
rect 24252 12448 24278 12474
rect 27150 12469 27176 12474
rect 27150 12452 27154 12469
rect 27154 12452 27171 12469
rect 27171 12452 27176 12469
rect 27150 12448 27176 12452
rect 25586 12435 25612 12440
rect 19146 12401 19172 12406
rect 19146 12384 19150 12401
rect 19150 12384 19167 12401
rect 19167 12384 19172 12401
rect 19146 12380 19172 12384
rect 18594 12346 18620 12372
rect 25586 12418 25588 12435
rect 25588 12418 25612 12435
rect 25586 12414 25612 12418
rect 27334 12435 27360 12440
rect 27334 12418 27338 12435
rect 27338 12418 27355 12435
rect 27355 12418 27360 12435
rect 27334 12414 27360 12418
rect 28116 12414 28142 12440
rect 28392 12414 28418 12440
rect 18318 12312 18344 12338
rect 19376 12312 19402 12338
rect 24436 12380 24462 12406
rect 25402 12380 25428 12406
rect 25632 12380 25658 12406
rect 26690 12380 26716 12406
rect 26782 12401 26808 12406
rect 26782 12384 26786 12401
rect 26786 12384 26803 12401
rect 26803 12384 26808 12401
rect 26782 12380 26808 12384
rect 26874 12380 26900 12406
rect 24068 12367 24094 12372
rect 24068 12350 24072 12367
rect 24072 12350 24089 12367
rect 24089 12350 24094 12367
rect 24068 12346 24094 12350
rect 27196 12401 27222 12406
rect 27196 12384 27200 12401
rect 27200 12384 27217 12401
rect 27217 12384 27222 12401
rect 27196 12380 27222 12384
rect 14224 12278 14250 12304
rect 14914 12278 14940 12304
rect 16294 12299 16320 12304
rect 16294 12282 16298 12299
rect 16298 12282 16315 12299
rect 16315 12282 16320 12299
rect 16294 12278 16320 12282
rect 16984 12278 17010 12304
rect 17536 12278 17562 12304
rect 18502 12278 18528 12304
rect 19422 12278 19448 12304
rect 21492 12278 21518 12304
rect 23930 12299 23956 12304
rect 23930 12282 23934 12299
rect 23934 12282 23951 12299
rect 23951 12282 23956 12299
rect 23930 12278 23956 12282
rect 26828 12278 26854 12304
rect 27380 12401 27406 12406
rect 27380 12384 27384 12401
rect 27384 12384 27401 12401
rect 27401 12384 27406 12401
rect 27380 12380 27406 12384
rect 29680 12380 29706 12406
rect 27840 12346 27866 12372
rect 28116 12367 28142 12372
rect 28116 12350 28120 12367
rect 28120 12350 28137 12367
rect 28137 12350 28142 12367
rect 28116 12346 28142 12350
rect 29588 12278 29614 12304
rect 7416 12197 7442 12202
rect 7416 12180 7420 12197
rect 7420 12180 7437 12197
rect 7437 12180 7442 12197
rect 7416 12176 7442 12180
rect 11556 12176 11582 12202
rect 13994 12176 14020 12202
rect 14684 12176 14710 12202
rect 15696 12176 15722 12202
rect 16800 12176 16826 12202
rect 19146 12176 19172 12202
rect 5392 12142 5418 12168
rect 4518 12108 4544 12134
rect 5852 12074 5878 12100
rect 5944 12095 5970 12100
rect 5944 12078 5965 12095
rect 5965 12078 5970 12095
rect 5944 12074 5970 12078
rect 4840 12061 4866 12066
rect 4840 12044 4844 12061
rect 4844 12044 4861 12061
rect 4861 12044 4866 12061
rect 4840 12040 4866 12044
rect 5530 12040 5556 12066
rect 5668 12040 5694 12066
rect 7324 12074 7350 12100
rect 7416 12095 7442 12100
rect 7416 12078 7420 12095
rect 7420 12078 7437 12095
rect 7437 12078 7442 12095
rect 7416 12074 7442 12078
rect 7462 12095 7488 12100
rect 7462 12078 7466 12095
rect 7466 12078 7483 12095
rect 7483 12078 7488 12095
rect 7462 12074 7488 12078
rect 7554 12095 7580 12100
rect 7554 12078 7558 12095
rect 7558 12078 7575 12095
rect 7575 12078 7580 12095
rect 7554 12074 7580 12078
rect 8474 12108 8500 12134
rect 10038 12108 10064 12134
rect 11970 12129 11996 12134
rect 11970 12112 11974 12129
rect 11974 12112 11991 12129
rect 11991 12112 11996 12129
rect 11970 12108 11996 12112
rect 13856 12108 13882 12134
rect 9118 12074 9144 12100
rect 10222 12074 10248 12100
rect 10452 12074 10478 12100
rect 12016 12095 12042 12100
rect 12016 12078 12023 12095
rect 12023 12078 12040 12095
rect 12040 12078 12042 12095
rect 12016 12074 12042 12078
rect 12798 12074 12824 12100
rect 14224 12095 14250 12100
rect 14224 12078 14228 12095
rect 14228 12078 14245 12095
rect 14245 12078 14250 12095
rect 14224 12074 14250 12078
rect 14408 12095 14434 12100
rect 14408 12078 14415 12095
rect 14415 12078 14432 12095
rect 14432 12078 14434 12095
rect 16110 12142 16136 12168
rect 14408 12074 14434 12078
rect 14822 12095 14848 12100
rect 14822 12078 14826 12095
rect 14826 12078 14843 12095
rect 14843 12078 14848 12095
rect 14822 12074 14848 12078
rect 14914 12095 14940 12100
rect 14914 12078 14918 12095
rect 14918 12078 14935 12095
rect 14935 12078 14940 12095
rect 14914 12074 14940 12078
rect 15926 12095 15952 12100
rect 15926 12078 15930 12095
rect 15930 12078 15947 12095
rect 15947 12078 15952 12095
rect 15926 12074 15952 12078
rect 16110 12074 16136 12100
rect 16984 12095 17010 12100
rect 16984 12078 16988 12095
rect 16988 12078 17005 12095
rect 17005 12078 17010 12095
rect 16984 12074 17010 12078
rect 8566 12040 8592 12066
rect 8796 12040 8822 12066
rect 10406 12061 10432 12066
rect 10406 12044 10408 12061
rect 10408 12044 10432 12061
rect 10406 12040 10432 12044
rect 11832 12061 11858 12066
rect 11832 12044 11836 12061
rect 11836 12044 11853 12061
rect 11853 12044 11858 12061
rect 11832 12040 11858 12044
rect 11924 12061 11950 12066
rect 11924 12044 11928 12061
rect 11928 12044 11945 12061
rect 11945 12044 11950 12061
rect 11924 12040 11950 12044
rect 11970 12061 11996 12066
rect 11970 12044 11974 12061
rect 11974 12044 11991 12061
rect 11991 12044 11996 12061
rect 11970 12040 11996 12044
rect 12890 12040 12916 12066
rect 13166 12061 13192 12066
rect 13166 12044 13168 12061
rect 13168 12044 13192 12061
rect 13166 12040 13192 12044
rect 9532 12006 9558 12032
rect 15788 12061 15814 12066
rect 15788 12044 15792 12061
rect 15792 12044 15809 12061
rect 15809 12044 15814 12061
rect 15788 12040 15814 12044
rect 16294 12040 16320 12066
rect 16570 12040 16596 12066
rect 17260 12074 17286 12100
rect 19284 12142 19310 12168
rect 19514 12163 19540 12168
rect 19514 12146 19518 12163
rect 19518 12146 19535 12163
rect 19535 12146 19540 12163
rect 19514 12142 19540 12146
rect 18502 12129 18528 12134
rect 18502 12112 18506 12129
rect 18506 12112 18523 12129
rect 18523 12112 18528 12129
rect 18502 12108 18528 12112
rect 18640 12108 18666 12134
rect 17536 12095 17562 12100
rect 17536 12078 17540 12095
rect 17540 12078 17557 12095
rect 17557 12078 17562 12095
rect 17536 12074 17562 12078
rect 17904 12074 17930 12100
rect 19882 12095 19908 12100
rect 19882 12078 19886 12095
rect 19886 12078 19903 12095
rect 19903 12078 19908 12095
rect 19882 12074 19908 12078
rect 19376 12040 19402 12066
rect 22596 12108 22622 12134
rect 25402 12176 25428 12202
rect 26782 12176 26808 12202
rect 22090 12095 22116 12100
rect 22090 12078 22094 12095
rect 22094 12078 22111 12095
rect 22111 12078 22116 12095
rect 22090 12074 22116 12078
rect 25632 12074 25658 12100
rect 16662 12006 16688 12032
rect 17168 12006 17194 12032
rect 19468 12027 19494 12032
rect 19468 12010 19472 12027
rect 19472 12010 19489 12027
rect 19489 12010 19494 12027
rect 21584 12040 21610 12066
rect 25494 12040 25520 12066
rect 19468 12006 19494 12010
rect 4840 11904 4866 11930
rect 5392 11925 5418 11930
rect 5392 11908 5396 11925
rect 5396 11908 5413 11925
rect 5413 11908 5418 11925
rect 5392 11904 5418 11908
rect 5438 11925 5464 11930
rect 5438 11908 5442 11925
rect 5442 11908 5459 11925
rect 5459 11908 5464 11925
rect 5438 11904 5464 11908
rect 7324 11870 7350 11896
rect 5898 11836 5924 11862
rect 7094 11836 7120 11862
rect 8612 11836 8638 11862
rect 8934 11857 8960 11862
rect 8934 11840 8938 11857
rect 8938 11840 8955 11857
rect 8955 11840 8960 11857
rect 8934 11836 8960 11840
rect 8980 11836 9006 11862
rect 9118 11857 9144 11862
rect 9118 11840 9122 11857
rect 9122 11840 9139 11857
rect 9139 11840 9144 11857
rect 9118 11836 9144 11840
rect 11694 11904 11720 11930
rect 15788 11904 15814 11930
rect 19376 11925 19402 11930
rect 19376 11908 19380 11925
rect 19380 11908 19397 11925
rect 19397 11908 19402 11925
rect 19376 11904 19402 11908
rect 27196 11904 27222 11930
rect 9716 11870 9742 11896
rect 9992 11870 10018 11896
rect 13028 11891 13054 11896
rect 9532 11836 9558 11862
rect 9578 11857 9604 11862
rect 9578 11840 9582 11857
rect 9582 11840 9599 11857
rect 9599 11840 9604 11857
rect 9578 11836 9604 11840
rect 9670 11857 9696 11862
rect 9670 11840 9674 11857
rect 9674 11840 9691 11857
rect 9691 11840 9696 11857
rect 9670 11836 9696 11840
rect 10222 11836 10248 11862
rect 13028 11874 13030 11891
rect 13030 11874 13054 11891
rect 13028 11870 13054 11874
rect 5346 11802 5372 11828
rect 5484 11823 5510 11828
rect 5484 11806 5488 11823
rect 5488 11806 5505 11823
rect 5505 11806 5510 11823
rect 5484 11802 5510 11806
rect 6864 11823 6890 11828
rect 6864 11806 6868 11823
rect 6868 11806 6885 11823
rect 6885 11806 6890 11823
rect 6864 11802 6890 11806
rect 9900 11802 9926 11828
rect 12798 11857 12824 11862
rect 10866 11802 10892 11828
rect 12798 11840 12802 11857
rect 12802 11840 12819 11857
rect 12819 11840 12824 11857
rect 12798 11836 12824 11840
rect 12936 11857 12962 11862
rect 12936 11840 12957 11857
rect 12957 11840 12962 11857
rect 12936 11836 12962 11840
rect 14316 11857 14342 11862
rect 14316 11840 14320 11857
rect 14320 11840 14337 11857
rect 14337 11840 14342 11857
rect 14316 11836 14342 11840
rect 14362 11836 14388 11862
rect 14500 11857 14526 11862
rect 14500 11840 14507 11857
rect 14507 11840 14524 11857
rect 14524 11840 14526 11857
rect 14500 11836 14526 11840
rect 15972 11836 15998 11862
rect 16386 11870 16412 11896
rect 16248 11857 16274 11862
rect 16248 11840 16252 11857
rect 16252 11840 16269 11857
rect 16269 11840 16274 11857
rect 16248 11836 16274 11840
rect 16340 11836 16366 11862
rect 16524 11836 16550 11862
rect 18732 11836 18758 11862
rect 12384 11823 12410 11828
rect 12384 11806 12388 11823
rect 12388 11806 12405 11823
rect 12405 11806 12410 11823
rect 12384 11802 12410 11806
rect 20112 11836 20138 11862
rect 20480 11836 20506 11862
rect 21446 11870 21472 11896
rect 25632 11870 25658 11896
rect 26184 11870 26210 11896
rect 20756 11836 20782 11862
rect 20848 11836 20874 11862
rect 21630 11857 21656 11862
rect 21630 11840 21634 11857
rect 21634 11840 21651 11857
rect 21651 11840 21656 11857
rect 21630 11836 21656 11840
rect 21676 11857 21702 11862
rect 21676 11840 21680 11857
rect 21680 11840 21697 11857
rect 21697 11840 21702 11857
rect 21676 11836 21702 11840
rect 21722 11857 21748 11862
rect 21722 11840 21729 11857
rect 21729 11840 21746 11857
rect 21746 11840 21748 11857
rect 21722 11836 21748 11840
rect 25402 11836 25428 11862
rect 20158 11802 20184 11828
rect 21584 11823 21610 11828
rect 21584 11806 21588 11823
rect 21588 11806 21605 11823
rect 21605 11806 21610 11823
rect 21584 11802 21610 11806
rect 10866 11734 10892 11760
rect 14040 11768 14066 11794
rect 13166 11734 13192 11760
rect 19928 11734 19954 11760
rect 21722 11734 21748 11760
rect 7416 11632 7442 11658
rect 9578 11632 9604 11658
rect 9716 11632 9742 11658
rect 11648 11632 11674 11658
rect 11970 11632 11996 11658
rect 13074 11632 13100 11658
rect 14316 11632 14342 11658
rect 18732 11632 18758 11658
rect 5898 11551 5924 11556
rect 5898 11534 5902 11551
rect 5902 11534 5919 11551
rect 5919 11534 5924 11551
rect 5898 11530 5924 11534
rect 5944 11530 5970 11556
rect 6174 11530 6200 11556
rect 8474 11564 8500 11590
rect 10176 11564 10202 11590
rect 7600 11551 7626 11556
rect 7600 11534 7604 11551
rect 7604 11534 7621 11551
rect 7621 11534 7626 11551
rect 7600 11530 7626 11534
rect 8704 11530 8730 11556
rect 6128 11517 6154 11522
rect 6128 11500 6130 11517
rect 6130 11500 6154 11517
rect 6128 11496 6154 11500
rect 7554 11517 7580 11522
rect 7554 11500 7558 11517
rect 7558 11500 7575 11517
rect 7575 11500 7580 11517
rect 7554 11496 7580 11500
rect 8612 11496 8638 11522
rect 9900 11530 9926 11556
rect 10452 11564 10478 11590
rect 10866 11530 10892 11556
rect 12798 11564 12824 11590
rect 16662 11564 16688 11590
rect 17444 11564 17470 11590
rect 21170 11564 21196 11590
rect 11096 11551 11122 11556
rect 11096 11534 11117 11551
rect 11117 11534 11122 11551
rect 11096 11530 11122 11534
rect 9946 11496 9972 11522
rect 12982 11530 13008 11556
rect 16340 11551 16366 11556
rect 16340 11534 16344 11551
rect 16344 11534 16361 11551
rect 16361 11534 16366 11551
rect 16340 11530 16366 11534
rect 16386 11551 16412 11556
rect 16386 11534 16390 11551
rect 16390 11534 16407 11551
rect 16407 11534 16412 11551
rect 16386 11530 16412 11534
rect 18640 11551 18666 11556
rect 18640 11534 18644 11551
rect 18644 11534 18661 11551
rect 18661 11534 18666 11551
rect 18640 11530 18666 11534
rect 18732 11551 18758 11556
rect 18732 11534 18736 11551
rect 18736 11534 18753 11551
rect 18753 11534 18758 11551
rect 18732 11530 18758 11534
rect 19468 11551 19494 11556
rect 19468 11534 19472 11551
rect 19472 11534 19489 11551
rect 19489 11534 19494 11551
rect 19468 11530 19494 11534
rect 19836 11530 19862 11556
rect 19928 11530 19954 11556
rect 12936 11496 12962 11522
rect 13166 11517 13192 11522
rect 13166 11500 13168 11517
rect 13168 11500 13192 11517
rect 13166 11496 13192 11500
rect 18548 11496 18574 11522
rect 10314 11483 10340 11488
rect 10314 11466 10318 11483
rect 10318 11466 10335 11483
rect 10335 11466 10340 11483
rect 10314 11462 10340 11466
rect 16110 11462 16136 11488
rect 7600 11360 7626 11386
rect 9670 11360 9696 11386
rect 21676 11360 21702 11386
rect 24436 11381 24462 11386
rect 24436 11364 24440 11381
rect 24440 11364 24457 11381
rect 24457 11364 24462 11381
rect 24436 11360 24462 11364
rect 4748 11347 4774 11352
rect 4748 11330 4750 11347
rect 4750 11330 4774 11347
rect 4748 11326 4774 11330
rect 5760 11326 5786 11352
rect 6174 11326 6200 11352
rect 6864 11326 6890 11352
rect 4518 11313 4544 11318
rect 4518 11296 4522 11313
rect 4522 11296 4539 11313
rect 4539 11296 4544 11313
rect 4518 11292 4544 11296
rect 6404 11292 6430 11318
rect 16156 11292 16182 11318
rect 16570 11292 16596 11318
rect 17122 11313 17148 11318
rect 17122 11296 17126 11313
rect 17126 11296 17143 11313
rect 17143 11296 17148 11313
rect 17122 11292 17148 11296
rect 17444 11313 17470 11318
rect 17444 11296 17448 11313
rect 17448 11296 17465 11313
rect 17465 11296 17470 11313
rect 17444 11292 17470 11296
rect 17536 11313 17562 11318
rect 17536 11296 17540 11313
rect 17540 11296 17557 11313
rect 17557 11296 17562 11313
rect 17536 11292 17562 11296
rect 18410 11292 18436 11318
rect 18594 11326 18620 11352
rect 20710 11347 20736 11352
rect 20710 11330 20712 11347
rect 20712 11330 20736 11347
rect 20710 11326 20736 11330
rect 28346 11347 28372 11352
rect 28346 11330 28348 11347
rect 28348 11330 28372 11347
rect 28346 11326 28372 11330
rect 18548 11313 18574 11318
rect 18548 11296 18552 11313
rect 18552 11296 18569 11313
rect 18569 11296 18574 11313
rect 18548 11292 18574 11296
rect 20112 11292 20138 11318
rect 24298 11292 24324 11318
rect 5622 11258 5648 11284
rect 5898 11258 5924 11284
rect 7554 11258 7580 11284
rect 17076 11279 17102 11284
rect 17076 11262 17080 11279
rect 17080 11262 17097 11279
rect 17097 11262 17102 11279
rect 17076 11258 17102 11262
rect 17214 11279 17240 11284
rect 17214 11262 17218 11279
rect 17218 11262 17235 11279
rect 17235 11262 17240 11279
rect 17214 11258 17240 11262
rect 16248 11224 16274 11250
rect 20158 11258 20184 11284
rect 24574 11313 24600 11318
rect 24574 11296 24578 11313
rect 24578 11296 24595 11313
rect 24595 11296 24600 11313
rect 24574 11292 24600 11296
rect 28392 11292 28418 11318
rect 28668 11292 28694 11318
rect 28714 11292 28740 11318
rect 28852 11292 28878 11318
rect 5530 11190 5556 11216
rect 16202 11211 16228 11216
rect 16202 11194 16206 11211
rect 16206 11194 16223 11211
rect 16223 11194 16228 11211
rect 16202 11190 16228 11194
rect 16340 11190 16366 11216
rect 18594 11190 18620 11216
rect 24758 11258 24784 11284
rect 28116 11279 28142 11284
rect 28116 11262 28120 11279
rect 28120 11262 28137 11279
rect 28137 11262 28142 11279
rect 28116 11258 28142 11262
rect 21170 11190 21196 11216
rect 29450 11211 29476 11216
rect 29450 11194 29454 11211
rect 29454 11194 29471 11211
rect 29471 11194 29476 11211
rect 29450 11190 29476 11194
rect 18732 11088 18758 11114
rect 24574 11088 24600 11114
rect 29082 11088 29108 11114
rect 7462 11054 7488 11080
rect 17030 11054 17056 11080
rect 17122 11054 17148 11080
rect 5346 11041 5372 11046
rect 5346 11024 5350 11041
rect 5350 11024 5367 11041
rect 5367 11024 5372 11041
rect 5346 11020 5372 11024
rect 11832 11020 11858 11046
rect 13948 11041 13974 11046
rect 13948 11024 13952 11041
rect 13952 11024 13969 11041
rect 13969 11024 13974 11041
rect 13948 11020 13974 11024
rect 16340 11041 16366 11046
rect 16340 11024 16344 11041
rect 16344 11024 16361 11041
rect 16361 11024 16366 11041
rect 16340 11020 16366 11024
rect 17214 11041 17240 11046
rect 17214 11024 17218 11041
rect 17218 11024 17235 11041
rect 17235 11024 17240 11041
rect 17214 11020 17240 11024
rect 5530 10986 5556 11012
rect 5622 11007 5648 11012
rect 5622 10990 5626 11007
rect 5626 10990 5643 11007
rect 5643 10990 5648 11007
rect 5622 10986 5648 10990
rect 5760 11007 5786 11012
rect 5760 10990 5781 11007
rect 5781 10990 5786 11007
rect 5760 10986 5786 10990
rect 6910 10986 6936 11012
rect 10038 10986 10064 11012
rect 10866 10986 10892 11012
rect 11096 10986 11122 11012
rect 12614 10986 12640 11012
rect 14500 10986 14526 11012
rect 16156 10986 16182 11012
rect 16248 11007 16274 11012
rect 16248 10990 16252 11007
rect 16252 10990 16269 11007
rect 16269 10990 16274 11007
rect 16248 10986 16274 10990
rect 16386 11007 16412 11012
rect 16386 10990 16390 11007
rect 16390 10990 16407 11007
rect 16407 10990 16412 11007
rect 16386 10986 16412 10990
rect 11050 10973 11076 10978
rect 11050 10956 11052 10973
rect 11052 10956 11076 10973
rect 11050 10952 11076 10956
rect 17168 11007 17194 11012
rect 17168 10990 17172 11007
rect 17172 10990 17189 11007
rect 17189 10990 17194 11007
rect 17168 10986 17194 10990
rect 21170 11020 21196 11046
rect 22090 11020 22116 11046
rect 22918 11020 22944 11046
rect 26690 11020 26716 11046
rect 17904 10986 17930 11012
rect 18594 11007 18620 11012
rect 18594 10990 18598 11007
rect 18598 10990 18615 11007
rect 18615 10990 18620 11007
rect 18594 10986 18620 10990
rect 22688 11007 22714 11012
rect 22688 10990 22695 11007
rect 22695 10990 22712 11007
rect 22712 10990 22714 11007
rect 22688 10986 22714 10990
rect 23148 11007 23174 11012
rect 23148 10990 23152 11007
rect 23152 10990 23169 11007
rect 23169 10990 23174 11007
rect 23148 10986 23174 10990
rect 23240 11007 23266 11012
rect 23240 10990 23244 11007
rect 23244 10990 23261 11007
rect 23261 10990 23266 11007
rect 23240 10986 23266 10990
rect 23976 11007 24002 11012
rect 23976 10990 23980 11007
rect 23980 10990 23997 11007
rect 23997 10990 24002 11007
rect 23976 10986 24002 10990
rect 17260 10952 17286 10978
rect 18318 10952 18344 10978
rect 21216 10952 21242 10978
rect 21446 10973 21472 10978
rect 21446 10956 21448 10973
rect 21448 10956 21472 10973
rect 21446 10952 21472 10956
rect 22596 10973 22622 10978
rect 22596 10956 22600 10973
rect 22600 10956 22617 10973
rect 22617 10956 22622 10973
rect 22596 10952 22622 10956
rect 22642 10973 22668 10978
rect 22642 10956 22646 10973
rect 22646 10956 22663 10973
rect 22663 10956 22668 10973
rect 22642 10952 22668 10956
rect 23010 10952 23036 10978
rect 5116 10918 5142 10944
rect 5208 10939 5234 10944
rect 5208 10922 5212 10939
rect 5212 10922 5229 10939
rect 5229 10922 5234 10939
rect 5208 10918 5234 10922
rect 13672 10939 13698 10944
rect 13672 10922 13676 10939
rect 13676 10922 13693 10939
rect 13693 10922 13698 10939
rect 13672 10918 13698 10922
rect 13856 10939 13882 10944
rect 13856 10922 13860 10939
rect 13860 10922 13877 10939
rect 13877 10922 13882 10939
rect 13856 10918 13882 10922
rect 13902 10939 13928 10944
rect 13902 10922 13906 10939
rect 13906 10922 13923 10939
rect 13923 10922 13928 10939
rect 13902 10918 13928 10922
rect 15880 10918 15906 10944
rect 23194 10939 23220 10944
rect 23194 10922 23198 10939
rect 23198 10922 23215 10939
rect 23215 10922 23220 10939
rect 23194 10918 23220 10922
rect 24022 10939 24048 10944
rect 24022 10922 24026 10939
rect 24026 10922 24043 10939
rect 24043 10922 24048 10939
rect 24022 10918 24048 10922
rect 4748 10782 4774 10808
rect 10038 10769 10064 10774
rect 10038 10752 10042 10769
rect 10042 10752 10059 10769
rect 10059 10752 10064 10769
rect 10038 10748 10064 10752
rect 10314 10748 10340 10774
rect 11878 10714 11904 10740
rect 13902 10816 13928 10842
rect 15742 10816 15768 10842
rect 16524 10816 16550 10842
rect 20342 10816 20368 10842
rect 22642 10816 22668 10842
rect 23240 10816 23266 10842
rect 23516 10816 23542 10842
rect 12430 10782 12456 10808
rect 12614 10803 12640 10808
rect 12614 10786 12616 10803
rect 12616 10786 12640 10803
rect 12614 10782 12640 10786
rect 14500 10782 14526 10808
rect 14730 10748 14756 10774
rect 15144 10748 15170 10774
rect 12384 10735 12410 10740
rect 12384 10718 12388 10735
rect 12388 10718 12405 10735
rect 12405 10718 12410 10735
rect 12384 10714 12410 10718
rect 14040 10714 14066 10740
rect 5346 10646 5372 10672
rect 10682 10646 10708 10672
rect 18732 10748 18758 10774
rect 17536 10714 17562 10740
rect 18318 10735 18344 10740
rect 18318 10718 18322 10735
rect 18322 10718 18339 10735
rect 18339 10718 18344 10735
rect 18318 10714 18344 10718
rect 18640 10646 18666 10672
rect 19928 10782 19954 10808
rect 20894 10782 20920 10808
rect 21354 10782 21380 10808
rect 23194 10782 23220 10808
rect 24022 10782 24048 10808
rect 26828 10837 26854 10842
rect 26828 10820 26832 10837
rect 26832 10820 26849 10837
rect 26849 10820 26854 10837
rect 26828 10816 26854 10820
rect 29082 10837 29108 10842
rect 29082 10820 29086 10837
rect 29086 10820 29103 10837
rect 29103 10820 29108 10837
rect 29082 10816 29108 10820
rect 25586 10803 25612 10808
rect 25586 10786 25588 10803
rect 25588 10786 25612 10803
rect 25586 10782 25612 10786
rect 29496 10782 29522 10808
rect 20296 10769 20322 10774
rect 20296 10752 20300 10769
rect 20300 10752 20317 10769
rect 20317 10752 20322 10769
rect 20296 10748 20322 10752
rect 20434 10748 20460 10774
rect 21216 10769 21242 10774
rect 20112 10714 20138 10740
rect 21216 10752 21237 10769
rect 21237 10752 21242 10769
rect 21216 10748 21242 10752
rect 22918 10769 22944 10774
rect 22918 10752 22922 10769
rect 22922 10752 22939 10769
rect 22939 10752 22944 10769
rect 22918 10748 22944 10752
rect 23102 10748 23128 10774
rect 19928 10680 19954 10706
rect 19330 10646 19356 10672
rect 20158 10646 20184 10672
rect 20618 10646 20644 10672
rect 23240 10735 23266 10740
rect 23240 10718 23244 10735
rect 23244 10718 23261 10735
rect 23261 10718 23266 10735
rect 23240 10714 23266 10718
rect 25678 10748 25704 10774
rect 27012 10748 27038 10774
rect 28944 10748 28970 10774
rect 29450 10748 29476 10774
rect 21170 10646 21196 10672
rect 23240 10646 23266 10672
rect 23562 10646 23588 10672
rect 24666 10714 24692 10740
rect 24804 10714 24830 10740
rect 25356 10735 25382 10740
rect 25356 10718 25360 10735
rect 25360 10718 25377 10735
rect 25377 10718 25382 10735
rect 25356 10714 25382 10718
rect 26230 10714 26256 10740
rect 24620 10646 24646 10672
rect 24896 10646 24922 10672
rect 25678 10646 25704 10672
rect 26276 10646 26302 10672
rect 26736 10667 26762 10672
rect 26736 10650 26740 10667
rect 26740 10650 26757 10667
rect 26757 10650 26762 10667
rect 26736 10646 26762 10650
rect 5622 10544 5648 10570
rect 5116 10497 5142 10502
rect 5116 10480 5120 10497
rect 5120 10480 5137 10497
rect 5137 10480 5142 10497
rect 5116 10476 5142 10480
rect 8474 10476 8500 10502
rect 5668 10442 5694 10468
rect 7600 10442 7626 10468
rect 8336 10463 8362 10468
rect 8336 10446 8340 10463
rect 8340 10446 8357 10463
rect 8357 10446 8362 10463
rect 8336 10442 8362 10446
rect 9256 10544 9282 10570
rect 10682 10544 10708 10570
rect 13948 10544 13974 10570
rect 17260 10544 17286 10570
rect 18732 10544 18758 10570
rect 20296 10544 20322 10570
rect 23010 10565 23036 10570
rect 23010 10548 23014 10565
rect 23014 10548 23031 10565
rect 23031 10548 23036 10565
rect 23010 10544 23036 10548
rect 23148 10544 23174 10570
rect 23976 10544 24002 10570
rect 24114 10544 24140 10570
rect 14776 10531 14802 10536
rect 14776 10514 14780 10531
rect 14780 10514 14797 10531
rect 14797 10514 14802 10531
rect 14776 10510 14802 10514
rect 20342 10510 20368 10536
rect 9532 10476 9558 10502
rect 13672 10497 13698 10502
rect 13672 10480 13676 10497
rect 13676 10480 13693 10497
rect 13693 10480 13698 10497
rect 13672 10476 13698 10480
rect 13856 10476 13882 10502
rect 13948 10476 13974 10502
rect 16202 10476 16228 10502
rect 19330 10476 19356 10502
rect 24620 10497 24646 10502
rect 24620 10480 24624 10497
rect 24624 10480 24641 10497
rect 24641 10480 24646 10497
rect 24620 10476 24646 10480
rect 12384 10442 12410 10468
rect 5208 10374 5234 10400
rect 9026 10408 9052 10434
rect 9578 10408 9604 10434
rect 8382 10395 8408 10400
rect 8382 10378 8386 10395
rect 8386 10378 8403 10395
rect 8403 10378 8408 10395
rect 8382 10374 8408 10378
rect 8934 10374 8960 10400
rect 9256 10374 9282 10400
rect 14408 10442 14434 10468
rect 15788 10442 15814 10468
rect 13902 10408 13928 10434
rect 14316 10408 14342 10434
rect 14592 10408 14618 10434
rect 17214 10463 17240 10468
rect 17214 10446 17218 10463
rect 17218 10446 17235 10463
rect 17235 10446 17240 10463
rect 17214 10442 17240 10446
rect 15972 10408 15998 10434
rect 16248 10408 16274 10434
rect 16524 10408 16550 10434
rect 18640 10463 18666 10468
rect 18640 10446 18644 10463
rect 18644 10446 18661 10463
rect 18661 10446 18666 10463
rect 18640 10442 18666 10446
rect 18686 10442 18712 10468
rect 20112 10442 20138 10468
rect 14040 10374 14066 10400
rect 14868 10395 14894 10400
rect 14868 10378 14872 10395
rect 14872 10378 14889 10395
rect 14889 10378 14894 10395
rect 14868 10374 14894 10378
rect 19652 10408 19678 10434
rect 17122 10374 17148 10400
rect 20020 10374 20046 10400
rect 23102 10463 23128 10468
rect 23102 10446 23106 10463
rect 23106 10446 23123 10463
rect 23123 10446 23128 10463
rect 23102 10442 23128 10446
rect 23516 10442 23542 10468
rect 24896 10442 24922 10468
rect 27610 10544 27636 10570
rect 28392 10544 28418 10570
rect 26690 10510 26716 10536
rect 26046 10463 26072 10468
rect 26046 10446 26063 10463
rect 26063 10446 26072 10463
rect 26276 10476 26302 10502
rect 26046 10442 26072 10446
rect 26230 10463 26256 10468
rect 26230 10446 26241 10463
rect 26241 10446 26256 10463
rect 26874 10476 26900 10502
rect 26230 10442 26256 10446
rect 27518 10463 27544 10468
rect 27518 10446 27522 10463
rect 27522 10446 27539 10463
rect 27539 10446 27544 10463
rect 27518 10442 27544 10446
rect 28944 10497 28970 10502
rect 28944 10480 28948 10497
rect 28948 10480 28965 10497
rect 28965 10480 28970 10497
rect 28944 10476 28970 10480
rect 28990 10463 29016 10468
rect 28990 10446 28997 10463
rect 28997 10446 29014 10463
rect 29014 10446 29016 10463
rect 28990 10442 29016 10446
rect 27564 10408 27590 10434
rect 27748 10429 27774 10434
rect 27748 10412 27750 10429
rect 27750 10412 27774 10429
rect 27748 10408 27774 10412
rect 29128 10408 29154 10434
rect 24160 10374 24186 10400
rect 24666 10374 24692 10400
rect 27150 10374 27176 10400
rect 7600 10272 7626 10298
rect 8152 10272 8178 10298
rect 9578 10272 9604 10298
rect 14316 10272 14342 10298
rect 9026 10259 9052 10264
rect 9026 10242 9030 10259
rect 9030 10242 9047 10259
rect 9047 10242 9052 10259
rect 9026 10238 9052 10242
rect 10544 10238 10570 10264
rect 14776 10238 14802 10264
rect 15880 10238 15906 10264
rect 22826 10272 22852 10298
rect 24114 10272 24140 10298
rect 26046 10272 26072 10298
rect 29128 10272 29154 10298
rect 16248 10238 16274 10264
rect 25586 10259 25612 10264
rect 25586 10242 25588 10259
rect 25588 10242 25612 10259
rect 25586 10238 25612 10242
rect 28346 10259 28372 10264
rect 28346 10242 28348 10259
rect 28348 10242 28372 10259
rect 28346 10238 28372 10242
rect 8382 10204 8408 10230
rect 8842 10225 8868 10230
rect 8842 10208 8846 10225
rect 8846 10208 8863 10225
rect 8863 10208 8868 10225
rect 8842 10204 8868 10208
rect 8934 10225 8960 10230
rect 8934 10208 8938 10225
rect 8938 10208 8955 10225
rect 8955 10208 8960 10225
rect 8934 10204 8960 10208
rect 9532 10225 9558 10230
rect 9532 10208 9536 10225
rect 9536 10208 9553 10225
rect 9553 10208 9558 10225
rect 9532 10204 9558 10208
rect 7508 10170 7534 10196
rect 9670 10191 9696 10196
rect 9670 10174 9674 10191
rect 9674 10174 9691 10191
rect 9691 10174 9696 10191
rect 9670 10170 9696 10174
rect 9716 10170 9742 10196
rect 14040 10170 14066 10196
rect 25356 10225 25382 10230
rect 25356 10208 25360 10225
rect 25360 10208 25377 10225
rect 25377 10208 25382 10225
rect 25356 10204 25382 10208
rect 25678 10204 25704 10230
rect 27610 10204 27636 10230
rect 27978 10204 28004 10230
rect 28116 10225 28142 10230
rect 28116 10208 28120 10225
rect 28120 10208 28137 10225
rect 28137 10208 28142 10225
rect 28116 10204 28142 10208
rect 28392 10204 28418 10230
rect 15972 10170 15998 10196
rect 17214 10170 17240 10196
rect 7922 10102 7948 10128
rect 14638 10102 14664 10128
rect 14868 10102 14894 10128
rect 7508 10021 7534 10026
rect 7508 10004 7512 10021
rect 7512 10004 7529 10021
rect 7529 10004 7534 10021
rect 7508 10000 7534 10004
rect 7922 9953 7948 9958
rect 7922 9936 7926 9953
rect 7926 9936 7943 9953
rect 7943 9936 7948 9953
rect 7922 9932 7948 9936
rect 8428 9932 8454 9958
rect 8888 9932 8914 9958
rect 7554 9919 7580 9924
rect 7554 9902 7558 9919
rect 7558 9902 7575 9919
rect 7575 9902 7580 9919
rect 7554 9898 7580 9902
rect 7600 9898 7626 9924
rect 8980 9898 9006 9924
rect 9256 9898 9282 9924
rect 9670 10021 9696 10026
rect 9670 10004 9674 10021
rect 9674 10004 9691 10021
rect 9691 10004 9696 10021
rect 9670 10000 9696 10004
rect 9532 9966 9558 9992
rect 9578 9953 9604 9958
rect 9578 9936 9582 9953
rect 9582 9936 9599 9953
rect 9599 9936 9604 9953
rect 9578 9932 9604 9936
rect 15972 9966 15998 9992
rect 9716 9898 9742 9924
rect 14408 9919 14434 9924
rect 14408 9902 14412 9919
rect 14412 9902 14429 9919
rect 14429 9902 14434 9919
rect 14408 9898 14434 9902
rect 15098 9932 15124 9958
rect 17904 9953 17930 9958
rect 17904 9936 17908 9953
rect 17908 9936 17925 9953
rect 17925 9936 17930 9953
rect 17904 9932 17930 9936
rect 18318 9932 18344 9958
rect 14638 9898 14664 9924
rect 17122 9919 17148 9924
rect 17122 9902 17126 9919
rect 17126 9902 17143 9919
rect 17143 9902 17148 9919
rect 17122 9898 17148 9902
rect 17214 9898 17240 9924
rect 17858 9919 17884 9924
rect 17858 9902 17862 9919
rect 17862 9902 17879 9919
rect 17879 9902 17884 9919
rect 17858 9898 17884 9902
rect 19054 9966 19080 9992
rect 23102 9966 23128 9992
rect 22642 9932 22668 9958
rect 19330 9898 19356 9924
rect 22688 9898 22714 9924
rect 7876 9864 7902 9890
rect 8152 9864 8178 9890
rect 9072 9851 9098 9856
rect 9072 9834 9076 9851
rect 9076 9834 9093 9851
rect 9093 9834 9098 9851
rect 9072 9830 9098 9834
rect 10314 9885 10340 9890
rect 10314 9868 10318 9885
rect 10318 9868 10335 9885
rect 10335 9868 10340 9885
rect 10314 9864 10340 9868
rect 10544 9864 10570 9890
rect 10820 9864 10846 9890
rect 13902 9864 13928 9890
rect 14592 9864 14618 9890
rect 9992 9830 10018 9856
rect 15236 9830 15262 9856
rect 22320 9885 22346 9890
rect 22320 9868 22324 9885
rect 22324 9868 22341 9885
rect 22341 9868 22346 9885
rect 22320 9864 22346 9868
rect 22550 9885 22576 9890
rect 22550 9868 22554 9885
rect 22554 9868 22571 9885
rect 22571 9868 22576 9885
rect 22550 9864 22576 9868
rect 22734 9864 22760 9890
rect 22182 9830 22208 9856
rect 27242 9830 27268 9856
rect 28484 9830 28510 9856
rect 28622 9830 28648 9856
rect 8888 9749 8914 9754
rect 8888 9732 8892 9749
rect 8892 9732 8909 9749
rect 8909 9732 8914 9749
rect 8888 9728 8914 9732
rect 7876 9694 7902 9720
rect 8106 9694 8132 9720
rect 8336 9694 8362 9720
rect 8934 9694 8960 9720
rect 7554 9660 7580 9686
rect 7876 9647 7902 9652
rect 7876 9630 7880 9647
rect 7880 9630 7897 9647
rect 7897 9630 7902 9647
rect 7876 9626 7902 9630
rect 14408 9728 14434 9754
rect 20618 9749 20644 9754
rect 20618 9732 20622 9749
rect 20622 9732 20639 9749
rect 20639 9732 20644 9749
rect 20618 9728 20644 9732
rect 23424 9749 23450 9754
rect 23424 9732 23428 9749
rect 23428 9732 23445 9749
rect 23445 9732 23450 9749
rect 23424 9728 23450 9732
rect 9716 9694 9742 9720
rect 15052 9694 15078 9720
rect 17030 9694 17056 9720
rect 17214 9694 17240 9720
rect 19238 9694 19264 9720
rect 9578 9681 9604 9686
rect 9578 9664 9582 9681
rect 9582 9664 9599 9681
rect 9599 9664 9604 9681
rect 9578 9660 9604 9664
rect 9992 9681 10018 9686
rect 9992 9664 9996 9681
rect 9996 9664 10013 9681
rect 10013 9664 10018 9681
rect 9992 9660 10018 9664
rect 14500 9681 14526 9686
rect 14500 9664 14504 9681
rect 14504 9664 14521 9681
rect 14521 9664 14526 9681
rect 14500 9660 14526 9664
rect 17122 9660 17148 9686
rect 19100 9681 19126 9686
rect 19100 9664 19104 9681
rect 19104 9664 19121 9681
rect 19121 9664 19126 9681
rect 19100 9660 19126 9664
rect 19146 9681 19172 9686
rect 19146 9664 19150 9681
rect 19150 9664 19167 9681
rect 19167 9664 19172 9681
rect 19146 9660 19172 9664
rect 22320 9694 22346 9720
rect 22642 9694 22668 9720
rect 20572 9681 20598 9686
rect 20572 9664 20576 9681
rect 20576 9664 20593 9681
rect 20593 9664 20598 9681
rect 20572 9660 20598 9664
rect 22550 9660 22576 9686
rect 22688 9681 22714 9686
rect 22688 9664 22692 9681
rect 22692 9664 22709 9681
rect 22709 9664 22714 9681
rect 22688 9660 22714 9664
rect 22734 9660 22760 9686
rect 25356 9694 25382 9720
rect 27242 9694 27268 9720
rect 28990 9694 29016 9720
rect 25632 9660 25658 9686
rect 8474 9626 8500 9652
rect 8888 9626 8914 9652
rect 10314 9626 10340 9652
rect 16570 9626 16596 9652
rect 16938 9626 16964 9652
rect 19008 9647 19034 9652
rect 19008 9630 19012 9647
rect 19012 9630 19029 9647
rect 19029 9630 19034 9647
rect 19008 9626 19034 9630
rect 8842 9613 8868 9618
rect 8842 9596 8846 9613
rect 8846 9596 8863 9613
rect 8863 9596 8868 9613
rect 8842 9592 8868 9596
rect 19882 9592 19908 9618
rect 22090 9626 22116 9652
rect 25356 9626 25382 9652
rect 28300 9626 28326 9652
rect 28438 9626 28464 9652
rect 29404 9626 29430 9652
rect 21722 9592 21748 9618
rect 24620 9592 24646 9618
rect 26966 9592 26992 9618
rect 28852 9592 28878 9618
rect 7784 9558 7810 9584
rect 14362 9579 14388 9584
rect 14362 9562 14366 9579
rect 14366 9562 14383 9579
rect 14383 9562 14388 9579
rect 14362 9558 14388 9562
rect 25862 9558 25888 9584
rect 28668 9558 28694 9584
rect 15052 9477 15078 9482
rect 15052 9460 15056 9477
rect 15056 9460 15073 9477
rect 15073 9460 15078 9477
rect 15052 9456 15078 9460
rect 20572 9456 20598 9482
rect 23976 9456 24002 9482
rect 26690 9456 26716 9482
rect 26736 9456 26762 9482
rect 21400 9422 21426 9448
rect 23884 9422 23910 9448
rect 7784 9409 7810 9414
rect 7784 9392 7788 9409
rect 7788 9392 7805 9409
rect 7805 9392 7810 9409
rect 7784 9388 7810 9392
rect 8888 9388 8914 9414
rect 7600 9354 7626 9380
rect 14040 9375 14066 9380
rect 14040 9358 14044 9375
rect 14044 9358 14061 9375
rect 14061 9358 14066 9375
rect 14040 9354 14066 9358
rect 14362 9354 14388 9380
rect 14408 9354 14434 9380
rect 15098 9409 15124 9414
rect 15098 9392 15102 9409
rect 15102 9392 15119 9409
rect 15119 9392 15124 9409
rect 15098 9388 15124 9392
rect 19008 9388 19034 9414
rect 7738 9320 7764 9346
rect 8152 9320 8178 9346
rect 14546 9286 14572 9312
rect 16110 9354 16136 9380
rect 18640 9354 18666 9380
rect 19100 9354 19126 9380
rect 19284 9354 19310 9380
rect 15466 9320 15492 9346
rect 19146 9320 19172 9346
rect 19606 9375 19632 9380
rect 19606 9358 19610 9375
rect 19610 9358 19627 9375
rect 19627 9358 19632 9375
rect 19606 9354 19632 9358
rect 20250 9354 20276 9380
rect 21354 9388 21380 9414
rect 20664 9375 20690 9380
rect 20664 9358 20668 9375
rect 20668 9358 20685 9375
rect 20685 9358 20690 9375
rect 20664 9354 20690 9358
rect 22182 9388 22208 9414
rect 22550 9388 22576 9414
rect 22780 9388 22806 9414
rect 23240 9388 23266 9414
rect 23838 9388 23864 9414
rect 25264 9409 25290 9414
rect 25264 9392 25268 9409
rect 25268 9392 25285 9409
rect 25285 9392 25290 9409
rect 25264 9388 25290 9392
rect 27058 9388 27084 9414
rect 27150 9409 27176 9414
rect 27150 9392 27154 9409
rect 27154 9392 27171 9409
rect 27171 9392 27176 9409
rect 27150 9388 27176 9392
rect 27978 9409 28004 9414
rect 27978 9392 27982 9409
rect 27982 9392 27999 9409
rect 27999 9392 28004 9409
rect 27978 9388 28004 9392
rect 20434 9320 20460 9346
rect 20526 9341 20552 9346
rect 20526 9324 20530 9341
rect 20530 9324 20547 9341
rect 20547 9324 20552 9341
rect 20526 9320 20552 9324
rect 21998 9320 22024 9346
rect 22642 9375 22668 9380
rect 22642 9358 22646 9375
rect 22646 9358 22663 9375
rect 22663 9358 22668 9375
rect 22642 9354 22668 9358
rect 22688 9354 22714 9380
rect 23424 9354 23450 9380
rect 26874 9354 26900 9380
rect 29036 9456 29062 9482
rect 29496 9477 29522 9482
rect 29496 9460 29500 9477
rect 29500 9460 29517 9477
rect 29517 9460 29522 9477
rect 29496 9456 29522 9460
rect 29174 9354 29200 9380
rect 29588 9375 29614 9380
rect 29588 9358 29592 9375
rect 29592 9358 29609 9375
rect 29609 9358 29614 9375
rect 29588 9354 29614 9358
rect 29680 9375 29706 9380
rect 29680 9358 29687 9375
rect 29687 9358 29704 9375
rect 29704 9358 29706 9375
rect 29680 9354 29706 9358
rect 15788 9307 15814 9312
rect 15788 9290 15792 9307
rect 15792 9290 15809 9307
rect 15809 9290 15814 9307
rect 15788 9286 15814 9290
rect 15880 9286 15906 9312
rect 18962 9286 18988 9312
rect 21952 9286 21978 9312
rect 22964 9307 22990 9312
rect 22964 9290 22968 9307
rect 22968 9290 22985 9307
rect 22985 9290 22990 9307
rect 22964 9286 22990 9290
rect 23976 9286 24002 9312
rect 24206 9341 24232 9346
rect 24206 9324 24208 9341
rect 24208 9324 24232 9341
rect 24206 9320 24232 9324
rect 25356 9341 25382 9346
rect 25356 9324 25360 9341
rect 25360 9324 25377 9341
rect 25377 9324 25382 9341
rect 25356 9320 25382 9324
rect 25402 9341 25428 9346
rect 25402 9324 25406 9341
rect 25406 9324 25423 9341
rect 25423 9324 25428 9341
rect 25402 9320 25428 9324
rect 28024 9320 28050 9346
rect 28208 9341 28234 9346
rect 28208 9324 28210 9341
rect 28210 9324 28234 9341
rect 28208 9320 28234 9324
rect 29634 9341 29660 9346
rect 29634 9324 29638 9341
rect 29638 9324 29655 9341
rect 29655 9324 29660 9341
rect 29634 9320 29660 9324
rect 26920 9286 26946 9312
rect 27150 9286 27176 9312
rect 14500 9184 14526 9210
rect 13810 9150 13836 9176
rect 14408 9150 14434 9176
rect 14132 9116 14158 9142
rect 14546 9137 14572 9142
rect 14546 9120 14550 9137
rect 14550 9120 14567 9137
rect 14567 9120 14572 9137
rect 14546 9116 14572 9120
rect 14638 9150 14664 9176
rect 15926 9150 15952 9176
rect 15972 9116 15998 9142
rect 19238 9184 19264 9210
rect 20526 9184 20552 9210
rect 22596 9184 22622 9210
rect 23424 9205 23450 9210
rect 23424 9188 23428 9205
rect 23428 9188 23445 9205
rect 23445 9188 23450 9205
rect 23424 9184 23450 9188
rect 25402 9184 25428 9210
rect 26920 9205 26946 9210
rect 26920 9188 26924 9205
rect 26924 9188 26941 9205
rect 26941 9188 26946 9205
rect 26920 9184 26946 9188
rect 29634 9184 29660 9210
rect 18640 9150 18666 9176
rect 20066 9171 20092 9176
rect 20066 9154 20068 9171
rect 20068 9154 20092 9171
rect 20066 9150 20092 9154
rect 19146 9116 19172 9142
rect 14546 9048 14572 9074
rect 15466 9103 15492 9108
rect 15466 9086 15470 9103
rect 15470 9086 15487 9103
rect 15487 9086 15492 9103
rect 15466 9082 15492 9086
rect 14454 9014 14480 9040
rect 17076 9103 17102 9108
rect 17076 9086 17080 9103
rect 17080 9086 17097 9103
rect 17097 9086 17102 9103
rect 17076 9082 17102 9086
rect 17122 9103 17148 9108
rect 17122 9086 17126 9103
rect 17126 9086 17143 9103
rect 17143 9086 17148 9103
rect 17122 9082 17148 9086
rect 17168 9082 17194 9108
rect 18916 9082 18942 9108
rect 19238 9137 19264 9142
rect 19238 9120 19242 9137
rect 19242 9120 19259 9137
rect 19259 9120 19264 9137
rect 19238 9116 19264 9120
rect 19606 9116 19632 9142
rect 20112 9116 20138 9142
rect 20572 9116 20598 9142
rect 16018 9014 16044 9040
rect 17168 9035 17194 9040
rect 17168 9018 17172 9035
rect 17172 9018 17189 9035
rect 17189 9018 17194 9035
rect 17168 9014 17194 9018
rect 19376 9082 19402 9108
rect 19698 9082 19724 9108
rect 19284 9048 19310 9074
rect 20480 9014 20506 9040
rect 21998 9116 22024 9142
rect 22734 9150 22760 9176
rect 23884 9150 23910 9176
rect 25678 9150 25704 9176
rect 25862 9171 25888 9176
rect 25862 9154 25864 9171
rect 25864 9154 25888 9171
rect 25862 9150 25888 9154
rect 26874 9150 26900 9176
rect 22642 9116 22668 9142
rect 22780 9116 22806 9142
rect 23516 9116 23542 9142
rect 23976 9137 24002 9142
rect 23976 9120 23997 9137
rect 23997 9120 24002 9137
rect 23976 9116 24002 9120
rect 26920 9137 26946 9142
rect 26920 9120 26924 9137
rect 26924 9120 26941 9137
rect 26941 9120 26946 9137
rect 26920 9116 26946 9120
rect 23838 9103 23864 9108
rect 23838 9086 23842 9103
rect 23842 9086 23859 9103
rect 23859 9086 23864 9103
rect 23838 9082 23864 9086
rect 25632 9103 25658 9108
rect 25632 9086 25636 9103
rect 25636 9086 25653 9103
rect 25653 9086 25658 9103
rect 25632 9082 25658 9086
rect 27058 9137 27084 9142
rect 28024 9150 28050 9176
rect 27058 9120 27082 9137
rect 27082 9120 27084 9137
rect 27058 9116 27084 9120
rect 27242 9137 27268 9142
rect 27242 9120 27253 9137
rect 27253 9120 27268 9137
rect 27242 9116 27268 9120
rect 27610 9116 27636 9142
rect 27978 9116 28004 9142
rect 28438 9116 28464 9142
rect 27748 9082 27774 9108
rect 22688 9048 22714 9074
rect 24206 9014 24232 9040
rect 25816 9014 25842 9040
rect 14454 8912 14480 8938
rect 15972 8933 15998 8938
rect 15972 8916 15976 8933
rect 15976 8916 15993 8933
rect 15993 8916 15998 8933
rect 15972 8912 15998 8916
rect 17858 8933 17884 8938
rect 17858 8916 17862 8933
rect 17862 8916 17879 8933
rect 17879 8916 17884 8933
rect 17858 8912 17884 8916
rect 19928 8912 19954 8938
rect 5990 8844 6016 8870
rect 6036 8865 6062 8870
rect 6036 8848 6040 8865
rect 6040 8848 6057 8865
rect 6057 8848 6062 8865
rect 6036 8844 6062 8848
rect 7692 8865 7718 8870
rect 7692 8848 7696 8865
rect 7696 8848 7713 8865
rect 7713 8848 7718 8865
rect 7692 8844 7718 8848
rect 14132 8899 14158 8904
rect 14132 8882 14136 8899
rect 14136 8882 14153 8899
rect 14153 8882 14158 8899
rect 14132 8878 14158 8882
rect 14408 8878 14434 8904
rect 20710 8912 20736 8938
rect 5622 8810 5648 8836
rect 6082 8810 6108 8836
rect 7876 8810 7902 8836
rect 9532 8844 9558 8870
rect 10360 8865 10386 8870
rect 10360 8848 10364 8865
rect 10364 8848 10381 8865
rect 10381 8848 10386 8865
rect 10360 8844 10386 8848
rect 11096 8844 11122 8870
rect 8106 8831 8132 8836
rect 8106 8814 8110 8831
rect 8110 8814 8127 8831
rect 8127 8814 8132 8831
rect 8106 8810 8132 8814
rect 22044 8878 22070 8904
rect 18226 8844 18252 8870
rect 19698 8865 19724 8870
rect 19698 8848 19702 8865
rect 19702 8848 19719 8865
rect 19719 8848 19724 8865
rect 19698 8844 19724 8848
rect 22642 8844 22668 8870
rect 7830 8776 7856 8802
rect 10636 8776 10662 8802
rect 10820 8776 10846 8802
rect 11004 8776 11030 8802
rect 14316 8810 14342 8836
rect 13626 8776 13652 8802
rect 13856 8776 13882 8802
rect 15098 8810 15124 8836
rect 15236 8776 15262 8802
rect 15696 8797 15722 8802
rect 15696 8780 15700 8797
rect 15700 8780 15717 8797
rect 15717 8780 15722 8797
rect 15696 8776 15722 8780
rect 15788 8831 15814 8836
rect 15788 8814 15792 8831
rect 15792 8814 15809 8831
rect 15809 8814 15814 8831
rect 15788 8810 15814 8814
rect 15834 8831 15860 8836
rect 15834 8814 15838 8831
rect 15838 8814 15855 8831
rect 15855 8814 15860 8831
rect 15834 8810 15860 8814
rect 17168 8810 17194 8836
rect 17996 8831 18022 8836
rect 17996 8814 18000 8831
rect 18000 8814 18017 8831
rect 18017 8814 18022 8831
rect 17996 8810 18022 8814
rect 20112 8810 20138 8836
rect 20250 8810 20276 8836
rect 20388 8810 20414 8836
rect 22182 8831 22208 8836
rect 22182 8814 22186 8831
rect 22186 8814 22203 8831
rect 22203 8814 22208 8831
rect 22182 8810 22208 8814
rect 16570 8776 16596 8802
rect 17076 8776 17102 8802
rect 19054 8776 19080 8802
rect 19928 8797 19954 8802
rect 19928 8780 19930 8797
rect 19930 8780 19954 8797
rect 19928 8776 19954 8780
rect 21998 8776 22024 8802
rect 22780 8810 22806 8836
rect 27610 8912 27636 8938
rect 27748 8912 27774 8938
rect 22596 8776 22622 8802
rect 22688 8776 22714 8802
rect 25678 8776 25704 8802
rect 28346 8810 28372 8836
rect 7646 8763 7672 8768
rect 7646 8746 7650 8763
rect 7650 8746 7667 8763
rect 7667 8746 7672 8763
rect 7646 8742 7672 8746
rect 7784 8742 7810 8768
rect 14040 8742 14066 8768
rect 18410 8742 18436 8768
rect 22734 8763 22760 8768
rect 22734 8746 22738 8763
rect 22738 8746 22755 8763
rect 22755 8746 22760 8763
rect 22734 8742 22760 8746
rect 23608 8742 23634 8768
rect 25586 8742 25612 8768
rect 7646 8640 7672 8666
rect 7922 8640 7948 8666
rect 9532 8661 9558 8666
rect 9532 8644 9536 8661
rect 9536 8644 9553 8661
rect 9553 8644 9558 8661
rect 9532 8640 9558 8644
rect 7830 8627 7856 8632
rect 7830 8610 7834 8627
rect 7834 8610 7851 8627
rect 7851 8610 7856 8627
rect 7830 8606 7856 8610
rect 8106 8606 8132 8632
rect 8842 8606 8868 8632
rect 7738 8572 7764 8598
rect 7876 8572 7902 8598
rect 8520 8572 8546 8598
rect 9486 8593 9512 8598
rect 9486 8576 9490 8593
rect 9490 8576 9507 8593
rect 9507 8576 9512 8593
rect 9486 8572 9512 8576
rect 10452 8593 10478 8598
rect 10452 8576 10456 8593
rect 10456 8576 10473 8593
rect 10473 8576 10478 8593
rect 10452 8572 10478 8576
rect 10636 8606 10662 8632
rect 18410 8661 18436 8666
rect 18410 8644 18414 8661
rect 18414 8644 18431 8661
rect 18431 8644 18436 8661
rect 18410 8640 18436 8644
rect 22872 8661 22898 8666
rect 22872 8644 22876 8661
rect 22876 8644 22893 8661
rect 22893 8644 22898 8661
rect 22872 8640 22898 8644
rect 27058 8640 27084 8666
rect 21538 8606 21564 8632
rect 23608 8606 23634 8632
rect 25724 8606 25750 8632
rect 28806 8627 28832 8632
rect 28806 8610 28810 8627
rect 28810 8610 28827 8627
rect 28827 8610 28832 8627
rect 28806 8606 28832 8610
rect 28990 8606 29016 8632
rect 11050 8572 11076 8598
rect 17076 8593 17102 8598
rect 17076 8576 17080 8593
rect 17080 8576 17097 8593
rect 17097 8576 17102 8593
rect 17076 8572 17102 8576
rect 17168 8593 17194 8598
rect 17168 8576 17172 8593
rect 17172 8576 17189 8593
rect 17189 8576 17194 8593
rect 17168 8572 17194 8576
rect 18226 8593 18252 8598
rect 18226 8576 18230 8593
rect 18230 8576 18247 8593
rect 18247 8576 18252 8593
rect 18226 8572 18252 8576
rect 19238 8572 19264 8598
rect 21262 8593 21288 8598
rect 21262 8576 21266 8593
rect 21266 8576 21283 8593
rect 21283 8576 21288 8593
rect 21262 8572 21288 8576
rect 21308 8572 21334 8598
rect 21630 8593 21656 8598
rect 21630 8576 21634 8593
rect 21634 8576 21651 8593
rect 21651 8576 21656 8593
rect 21630 8572 21656 8576
rect 22182 8572 22208 8598
rect 22228 8572 22254 8598
rect 22596 8593 22622 8598
rect 22596 8576 22600 8593
rect 22600 8576 22617 8593
rect 22617 8576 22622 8593
rect 22596 8572 22622 8576
rect 22642 8572 22668 8598
rect 22780 8572 22806 8598
rect 23240 8572 23266 8598
rect 23516 8593 23542 8598
rect 23516 8576 23537 8593
rect 23537 8576 23542 8593
rect 23516 8572 23542 8576
rect 25678 8572 25704 8598
rect 28392 8572 28418 8598
rect 6358 8538 6384 8564
rect 6542 8559 6568 8564
rect 6542 8542 6546 8559
rect 6546 8542 6563 8559
rect 6563 8542 6568 8559
rect 6542 8538 6568 8542
rect 7692 8538 7718 8564
rect 9118 8538 9144 8564
rect 7876 8504 7902 8530
rect 8888 8504 8914 8530
rect 8980 8491 9006 8496
rect 8980 8474 8984 8491
rect 8984 8474 9001 8491
rect 9001 8474 9006 8491
rect 8980 8470 9006 8474
rect 10636 8559 10662 8564
rect 10636 8542 10640 8559
rect 10640 8542 10657 8559
rect 10657 8542 10662 8559
rect 10636 8538 10662 8542
rect 18272 8559 18298 8564
rect 18272 8542 18276 8559
rect 18276 8542 18293 8559
rect 18293 8542 18298 8559
rect 18272 8538 18298 8542
rect 22964 8559 22990 8564
rect 22964 8542 22968 8559
rect 22968 8542 22985 8559
rect 22985 8542 22990 8559
rect 22964 8538 22990 8542
rect 25816 8559 25842 8564
rect 25816 8542 25820 8559
rect 25820 8542 25837 8559
rect 25837 8542 25842 8559
rect 25816 8538 25842 8542
rect 28898 8593 28924 8598
rect 28898 8576 28905 8593
rect 28905 8576 28922 8593
rect 28922 8576 28924 8593
rect 28898 8572 28924 8576
rect 29128 8538 29154 8564
rect 17122 8504 17148 8530
rect 22136 8504 22162 8530
rect 22688 8504 22714 8530
rect 27150 8504 27176 8530
rect 11096 8470 11122 8496
rect 24344 8470 24370 8496
rect 8520 8389 8546 8394
rect 8520 8372 8524 8389
rect 8524 8372 8541 8389
rect 8541 8372 8546 8389
rect 8520 8368 8546 8372
rect 9486 8368 9512 8394
rect 19238 8334 19264 8360
rect 20342 8334 20368 8360
rect 21262 8334 21288 8360
rect 24298 8334 24324 8360
rect 24482 8368 24508 8394
rect 6036 8300 6062 8326
rect 6082 8300 6108 8326
rect 7784 8321 7810 8326
rect 7784 8304 7788 8321
rect 7788 8304 7805 8321
rect 7805 8304 7810 8321
rect 7784 8300 7810 8304
rect 20020 8300 20046 8326
rect 20388 8300 20414 8326
rect 7600 8266 7626 8292
rect 9532 8266 9558 8292
rect 19606 8287 19632 8292
rect 19606 8270 19610 8287
rect 19610 8270 19627 8287
rect 19627 8270 19632 8287
rect 19606 8266 19632 8270
rect 19790 8287 19816 8292
rect 19790 8270 19794 8287
rect 19794 8270 19811 8287
rect 19811 8270 19816 8287
rect 19790 8266 19816 8270
rect 6082 8232 6108 8258
rect 8750 8232 8776 8258
rect 19100 8232 19126 8258
rect 20894 8266 20920 8292
rect 21308 8266 21334 8292
rect 21998 8266 22024 8292
rect 22228 8287 22254 8292
rect 22228 8270 22232 8287
rect 22232 8270 22249 8287
rect 22249 8270 22254 8287
rect 22228 8266 22254 8270
rect 22642 8300 22668 8326
rect 22688 8266 22714 8292
rect 22780 8266 22806 8292
rect 22964 8266 22990 8292
rect 24344 8287 24370 8292
rect 24344 8270 24350 8287
rect 24350 8270 24370 8287
rect 24344 8266 24370 8270
rect 24390 8285 24416 8289
rect 24390 8268 24407 8285
rect 24407 8268 24416 8285
rect 24390 8263 24416 8268
rect 24513 8285 24539 8289
rect 24513 8268 24517 8285
rect 24517 8268 24534 8285
rect 24534 8268 24539 8285
rect 24513 8263 24539 8268
rect 24620 8266 24646 8292
rect 29358 8266 29384 8292
rect 6358 8198 6384 8224
rect 6864 8198 6890 8224
rect 7876 8198 7902 8224
rect 8842 8219 8868 8224
rect 8842 8202 8846 8219
rect 8846 8202 8863 8219
rect 8863 8202 8868 8219
rect 8842 8198 8868 8202
rect 20204 8198 20230 8224
rect 22918 8232 22944 8258
rect 26828 8232 26854 8258
rect 27380 8232 27406 8258
rect 22826 8198 22852 8224
rect 22964 8219 22990 8224
rect 22964 8202 22968 8219
rect 22968 8202 22985 8219
rect 22985 8202 22990 8219
rect 22964 8198 22990 8202
rect 23010 8198 23036 8224
rect 24298 8198 24324 8224
rect 24482 8219 24508 8224
rect 24482 8202 24486 8219
rect 24486 8202 24503 8219
rect 24503 8202 24508 8219
rect 24482 8198 24508 8202
rect 5990 8028 6016 8054
rect 6588 8028 6614 8054
rect 7692 8096 7718 8122
rect 7876 8096 7902 8122
rect 15696 8096 15722 8122
rect 17996 8096 18022 8122
rect 18272 8096 18298 8122
rect 19284 8096 19310 8122
rect 7738 8062 7764 8088
rect 7830 8062 7856 8088
rect 8198 8049 8224 8054
rect 8198 8032 8202 8049
rect 8202 8032 8219 8049
rect 8219 8032 8224 8049
rect 8198 8028 8224 8032
rect 20204 8062 20230 8088
rect 10452 8028 10478 8054
rect 10590 8028 10616 8054
rect 14408 8049 14434 8054
rect 14408 8032 14412 8049
rect 14412 8032 14429 8049
rect 14429 8032 14434 8049
rect 14408 8028 14434 8032
rect 14500 8049 14526 8054
rect 14500 8032 14504 8049
rect 14504 8032 14521 8049
rect 14521 8032 14526 8049
rect 14500 8028 14526 8032
rect 14546 8049 14572 8054
rect 14546 8032 14550 8049
rect 14550 8032 14567 8049
rect 14567 8032 14572 8049
rect 14546 8028 14572 8032
rect 16110 8028 16136 8054
rect 17490 8028 17516 8054
rect 18088 8028 18114 8054
rect 18640 8028 18666 8054
rect 6864 8015 6890 8020
rect 6864 7998 6868 8015
rect 6868 7998 6885 8015
rect 6885 7998 6890 8015
rect 6864 7994 6890 7998
rect 7646 7994 7672 8020
rect 7692 7994 7718 8020
rect 7922 7994 7948 8020
rect 10406 7994 10432 8020
rect 10636 7994 10662 8020
rect 13856 7994 13882 8020
rect 15880 7994 15906 8020
rect 15972 7994 15998 8020
rect 17398 8015 17424 8020
rect 17398 7998 17402 8015
rect 17402 7998 17419 8015
rect 17419 7998 17424 8015
rect 17398 7994 17424 7998
rect 19330 7994 19356 8020
rect 6818 7926 6844 7952
rect 8198 7960 8224 7986
rect 11556 7960 11582 7986
rect 17168 7960 17194 7986
rect 20342 8049 20368 8054
rect 20342 8032 20346 8049
rect 20346 8032 20363 8049
rect 20363 8032 20368 8049
rect 20342 8028 20368 8032
rect 20434 8083 20460 8088
rect 20434 8066 20438 8083
rect 20438 8066 20455 8083
rect 20455 8066 20460 8083
rect 21032 8096 21058 8122
rect 20434 8062 20460 8066
rect 20756 8028 20782 8054
rect 21078 8049 21104 8054
rect 21078 8032 21082 8049
rect 21082 8032 21099 8049
rect 21099 8032 21104 8049
rect 21078 8028 21104 8032
rect 21308 8096 21334 8122
rect 21354 8117 21380 8122
rect 21354 8100 21358 8117
rect 21358 8100 21375 8117
rect 21375 8100 21380 8117
rect 21354 8096 21380 8100
rect 22734 8096 22760 8122
rect 23010 8096 23036 8122
rect 24390 8096 24416 8122
rect 24482 8096 24508 8122
rect 24804 8117 24830 8122
rect 24804 8100 24808 8117
rect 24808 8100 24825 8117
rect 24825 8100 24830 8117
rect 24804 8096 24830 8100
rect 29128 8096 29154 8122
rect 23424 8083 23450 8088
rect 23424 8066 23426 8083
rect 23426 8066 23450 8083
rect 23424 8062 23450 8066
rect 28346 8083 28372 8088
rect 28346 8066 28348 8083
rect 28348 8066 28372 8083
rect 28346 8062 28372 8066
rect 21630 8028 21656 8054
rect 23240 8028 23266 8054
rect 23516 8028 23542 8054
rect 24712 8049 24738 8054
rect 24712 8032 24716 8049
rect 24716 8032 24733 8049
rect 24733 8032 24738 8049
rect 24712 8028 24738 8032
rect 25264 8028 25290 8054
rect 28070 8028 28096 8054
rect 28392 8028 28418 8054
rect 22136 7994 22162 8020
rect 22274 7994 22300 8020
rect 27978 7994 28004 8020
rect 20986 7960 21012 7986
rect 24758 7981 24784 7986
rect 24758 7964 24762 7981
rect 24762 7964 24779 7981
rect 24779 7964 24784 7981
rect 24758 7960 24784 7964
rect 7692 7926 7718 7952
rect 8106 7947 8132 7952
rect 8106 7930 8110 7947
rect 8110 7930 8127 7947
rect 8127 7930 8132 7947
rect 8106 7926 8132 7930
rect 10682 7926 10708 7952
rect 13718 7926 13744 7952
rect 20756 7926 20782 7952
rect 22136 7926 22162 7952
rect 22228 7926 22254 7952
rect 6542 7824 6568 7850
rect 8106 7824 8132 7850
rect 15972 7845 15998 7850
rect 15972 7828 15976 7845
rect 15976 7828 15993 7845
rect 15993 7828 15998 7845
rect 15972 7824 15998 7828
rect 17490 7845 17516 7850
rect 17490 7828 17494 7845
rect 17494 7828 17511 7845
rect 17511 7828 17516 7845
rect 17490 7824 17516 7828
rect 19652 7824 19678 7850
rect 28346 7824 28372 7850
rect 28990 7824 29016 7850
rect 29036 7824 29062 7850
rect 7646 7811 7672 7816
rect 7646 7794 7650 7811
rect 7650 7794 7667 7811
rect 7667 7794 7672 7811
rect 7646 7790 7672 7794
rect 14500 7790 14526 7816
rect 6588 7756 6614 7782
rect 6818 7743 6844 7748
rect 6818 7726 6822 7743
rect 6822 7726 6839 7743
rect 6839 7726 6844 7743
rect 6818 7722 6844 7726
rect 7784 7756 7810 7782
rect 10360 7756 10386 7782
rect 10682 7777 10708 7782
rect 10682 7760 10686 7777
rect 10686 7760 10703 7777
rect 10703 7760 10708 7777
rect 10682 7756 10708 7760
rect 7692 7722 7718 7748
rect 10406 7722 10432 7748
rect 13718 7743 13744 7748
rect 13718 7726 13722 7743
rect 13722 7726 13739 7743
rect 13739 7726 13744 7743
rect 13718 7722 13744 7726
rect 14040 7756 14066 7782
rect 13856 7743 13882 7748
rect 13856 7726 13860 7743
rect 13860 7726 13877 7743
rect 13877 7726 13882 7743
rect 13856 7722 13882 7726
rect 7922 7688 7948 7714
rect 11004 7688 11030 7714
rect 11510 7688 11536 7714
rect 14546 7722 14572 7748
rect 15972 7722 15998 7748
rect 19284 7790 19310 7816
rect 20020 7790 20046 7816
rect 20204 7790 20230 7816
rect 18272 7756 18298 7782
rect 18318 7722 18344 7748
rect 19146 7722 19172 7748
rect 20940 7756 20966 7782
rect 20020 7722 20046 7748
rect 22274 7790 22300 7816
rect 21538 7777 21564 7782
rect 21538 7760 21542 7777
rect 21542 7760 21559 7777
rect 21559 7760 21564 7777
rect 21538 7756 21564 7760
rect 21630 7756 21656 7782
rect 14408 7688 14434 7714
rect 19100 7688 19126 7714
rect 21446 7743 21472 7748
rect 21446 7726 21450 7743
rect 21450 7726 21467 7743
rect 21467 7726 21472 7743
rect 21446 7722 21472 7726
rect 22136 7722 22162 7748
rect 22182 7743 22208 7748
rect 22182 7726 22186 7743
rect 22186 7726 22203 7743
rect 22203 7726 22208 7743
rect 22182 7722 22208 7726
rect 22780 7756 22806 7782
rect 24804 7790 24830 7816
rect 22688 7722 22714 7748
rect 21078 7688 21104 7714
rect 26736 7743 26762 7748
rect 26736 7726 26740 7743
rect 26740 7726 26757 7743
rect 26757 7726 26762 7743
rect 26736 7722 26762 7726
rect 26828 7743 26854 7748
rect 26828 7726 26834 7743
rect 26834 7726 26854 7743
rect 26828 7722 26854 7726
rect 7830 7654 7856 7680
rect 8198 7654 8224 7680
rect 8750 7675 8776 7680
rect 8750 7658 8754 7675
rect 8754 7658 8771 7675
rect 8771 7658 8776 7675
rect 8750 7654 8776 7658
rect 19928 7675 19954 7680
rect 19928 7658 19932 7675
rect 19932 7658 19949 7675
rect 19949 7658 19954 7675
rect 19928 7654 19954 7658
rect 21676 7654 21702 7680
rect 24344 7654 24370 7680
rect 26874 7688 26900 7714
rect 27104 7722 27130 7748
rect 27978 7722 28004 7748
rect 28070 7743 28096 7748
rect 28070 7726 28091 7743
rect 28091 7726 28096 7743
rect 28070 7722 28096 7726
rect 27748 7688 27774 7714
rect 27886 7688 27912 7714
rect 28622 7722 28648 7748
rect 29312 7722 29338 7748
rect 29542 7743 29568 7748
rect 29542 7726 29546 7743
rect 29546 7726 29563 7743
rect 29563 7726 29568 7743
rect 29542 7722 29568 7726
rect 29726 7743 29752 7748
rect 29726 7726 29730 7743
rect 29730 7726 29747 7743
rect 29747 7726 29752 7743
rect 29726 7722 29752 7726
rect 29404 7688 29430 7714
rect 29680 7709 29706 7714
rect 29680 7692 29684 7709
rect 29684 7692 29701 7709
rect 29701 7692 29706 7709
rect 29680 7688 29706 7692
rect 27288 7654 27314 7680
rect 6174 7552 6200 7578
rect 15788 7552 15814 7578
rect 18272 7573 18298 7578
rect 18272 7556 18276 7573
rect 18276 7556 18293 7573
rect 18293 7556 18298 7573
rect 18272 7552 18298 7556
rect 5990 7518 6016 7544
rect 6082 7518 6108 7544
rect 7140 7539 7166 7544
rect 7140 7522 7144 7539
rect 7144 7522 7161 7539
rect 7161 7522 7166 7539
rect 7140 7518 7166 7522
rect 7692 7518 7718 7544
rect 11648 7539 11674 7544
rect 6220 7484 6246 7510
rect 7646 7484 7672 7510
rect 9072 7484 9098 7510
rect 9256 7505 9282 7510
rect 9256 7488 9260 7505
rect 9260 7488 9277 7505
rect 9277 7488 9282 7505
rect 9256 7484 9282 7488
rect 9440 7484 9466 7510
rect 9578 7484 9604 7510
rect 10406 7505 10432 7510
rect 10406 7488 10410 7505
rect 10410 7488 10427 7505
rect 10427 7488 10432 7505
rect 10406 7484 10432 7488
rect 11648 7522 11652 7539
rect 11652 7522 11669 7539
rect 11669 7522 11674 7539
rect 11648 7518 11674 7522
rect 19652 7518 19678 7544
rect 11096 7484 11122 7510
rect 11510 7484 11536 7510
rect 11832 7484 11858 7510
rect 15742 7484 15768 7510
rect 14316 7450 14342 7476
rect 18318 7505 18344 7510
rect 18318 7488 18322 7505
rect 18322 7488 18339 7505
rect 18339 7488 18344 7505
rect 18318 7484 18344 7488
rect 18962 7505 18988 7510
rect 18962 7488 18966 7505
rect 18966 7488 18983 7505
rect 18983 7488 18988 7505
rect 18962 7484 18988 7488
rect 19100 7505 19126 7510
rect 19100 7488 19104 7505
rect 19104 7488 19121 7505
rect 19121 7488 19126 7505
rect 19100 7484 19126 7488
rect 19330 7484 19356 7510
rect 20342 7484 20368 7510
rect 21446 7552 21472 7578
rect 24482 7552 24508 7578
rect 26874 7552 26900 7578
rect 29542 7552 29568 7578
rect 8198 7416 8224 7442
rect 9118 7416 9144 7442
rect 10590 7416 10616 7442
rect 6128 7382 6154 7408
rect 6588 7382 6614 7408
rect 6864 7382 6890 7408
rect 7600 7382 7626 7408
rect 7738 7382 7764 7408
rect 10406 7403 10432 7408
rect 10406 7386 10410 7403
rect 10410 7386 10427 7403
rect 10427 7386 10432 7403
rect 10406 7382 10432 7386
rect 10728 7403 10754 7408
rect 10728 7386 10732 7403
rect 10732 7386 10749 7403
rect 10749 7386 10754 7403
rect 10728 7382 10754 7386
rect 11556 7437 11582 7442
rect 11556 7420 11560 7437
rect 11560 7420 11577 7437
rect 11577 7420 11582 7437
rect 11556 7416 11582 7420
rect 20756 7539 20782 7544
rect 20756 7522 20760 7539
rect 20760 7522 20777 7539
rect 20777 7522 20782 7539
rect 20756 7518 20782 7522
rect 21032 7539 21058 7544
rect 21032 7522 21036 7539
rect 21036 7522 21053 7539
rect 21053 7522 21058 7539
rect 21032 7518 21058 7522
rect 21078 7539 21104 7544
rect 21078 7522 21082 7539
rect 21082 7522 21099 7539
rect 21099 7522 21104 7539
rect 21078 7518 21104 7522
rect 20986 7505 21012 7510
rect 20986 7488 20990 7505
rect 20990 7488 21007 7505
rect 21007 7488 21012 7505
rect 20986 7484 21012 7488
rect 22688 7450 22714 7476
rect 21400 7416 21426 7442
rect 20710 7382 20736 7408
rect 23516 7518 23542 7544
rect 25862 7518 25888 7544
rect 26092 7518 26118 7544
rect 28346 7539 28372 7544
rect 28346 7522 28348 7539
rect 28348 7522 28372 7539
rect 28346 7518 28372 7522
rect 23240 7484 23266 7510
rect 23562 7484 23588 7510
rect 26138 7484 26164 7510
rect 27978 7484 28004 7510
rect 28392 7484 28418 7510
rect 25816 7471 25842 7476
rect 25816 7454 25820 7471
rect 25820 7454 25837 7471
rect 25837 7454 25842 7471
rect 25816 7450 25842 7454
rect 23516 7382 23542 7408
rect 24666 7382 24692 7408
rect 8796 7280 8822 7306
rect 9072 7301 9098 7306
rect 9072 7284 9076 7301
rect 9076 7284 9093 7301
rect 9093 7284 9098 7301
rect 9072 7280 9098 7284
rect 10406 7280 10432 7306
rect 14316 7301 14342 7306
rect 14316 7284 14320 7301
rect 14320 7284 14337 7301
rect 14337 7284 14342 7301
rect 14316 7280 14342 7284
rect 21078 7280 21104 7306
rect 23240 7280 23266 7306
rect 25678 7280 25704 7306
rect 25816 7280 25842 7306
rect 6174 7212 6200 7238
rect 7600 7233 7626 7238
rect 7600 7216 7604 7233
rect 7604 7216 7621 7233
rect 7621 7216 7626 7233
rect 7600 7212 7626 7216
rect 7738 7233 7764 7238
rect 7738 7216 7742 7233
rect 7742 7216 7759 7233
rect 7759 7216 7764 7233
rect 7738 7212 7764 7216
rect 8106 7212 8132 7238
rect 5530 7199 5556 7204
rect 5530 7182 5534 7199
rect 5534 7182 5551 7199
rect 5551 7182 5556 7199
rect 5530 7178 5556 7182
rect 10590 7246 10616 7272
rect 11832 7246 11858 7272
rect 9026 7212 9052 7238
rect 10360 7212 10386 7238
rect 10820 7212 10846 7238
rect 11648 7233 11674 7238
rect 11648 7216 11652 7233
rect 11652 7216 11669 7233
rect 11669 7216 11674 7233
rect 11648 7212 11674 7216
rect 14040 7212 14066 7238
rect 5668 7165 5694 7170
rect 5668 7148 5672 7165
rect 5672 7148 5689 7165
rect 5689 7148 5694 7165
rect 5668 7144 5694 7148
rect 5944 7144 5970 7170
rect 6036 7144 6062 7170
rect 7600 7144 7626 7170
rect 7692 7144 7718 7170
rect 8888 7144 8914 7170
rect 9578 7199 9604 7204
rect 9578 7182 9582 7199
rect 9582 7182 9599 7199
rect 9599 7182 9604 7199
rect 9578 7178 9604 7182
rect 9440 7144 9466 7170
rect 11510 7178 11536 7204
rect 14408 7178 14434 7204
rect 15788 7178 15814 7204
rect 18640 7178 18666 7204
rect 18962 7212 18988 7238
rect 21400 7246 21426 7272
rect 19146 7212 19172 7238
rect 20066 7212 20092 7238
rect 22182 7212 22208 7238
rect 27748 7280 27774 7306
rect 27978 7246 28004 7272
rect 11004 7144 11030 7170
rect 18318 7144 18344 7170
rect 19606 7178 19632 7204
rect 19790 7178 19816 7204
rect 19974 7178 20000 7204
rect 22136 7178 22162 7204
rect 22642 7199 22668 7204
rect 22642 7182 22646 7199
rect 22646 7182 22663 7199
rect 22663 7182 22668 7199
rect 22642 7178 22668 7182
rect 22780 7178 22806 7204
rect 26138 7178 26164 7204
rect 20342 7144 20368 7170
rect 9302 7110 9328 7136
rect 11142 7110 11168 7136
rect 18410 7110 18436 7136
rect 19376 7110 19402 7136
rect 21308 7144 21334 7170
rect 24206 7144 24232 7170
rect 26966 7165 26992 7170
rect 26966 7148 26968 7165
rect 26968 7148 26992 7165
rect 26966 7144 26992 7148
rect 21124 7110 21150 7136
rect 21216 7110 21242 7136
rect 21446 7110 21472 7136
rect 22596 7110 22622 7136
rect 22918 7110 22944 7136
rect 24896 7110 24922 7136
rect 5668 7008 5694 7034
rect 8796 7008 8822 7034
rect 10728 7008 10754 7034
rect 10452 6974 10478 7000
rect 21124 7008 21150 7034
rect 13810 6995 13836 7000
rect 13810 6978 13814 6995
rect 13814 6978 13831 6995
rect 13831 6978 13836 6995
rect 13810 6974 13836 6978
rect 6128 6961 6154 6966
rect 6128 6944 6132 6961
rect 6132 6944 6149 6961
rect 6149 6944 6154 6961
rect 6128 6940 6154 6944
rect 8106 6940 8132 6966
rect 8888 6940 8914 6966
rect 11832 6940 11858 6966
rect 14270 6940 14296 6966
rect 15742 6974 15768 7000
rect 15788 6961 15814 6966
rect 6128 6872 6154 6898
rect 8198 6893 8224 6898
rect 8198 6876 8202 6893
rect 8202 6876 8219 6893
rect 8219 6876 8224 6893
rect 8198 6872 8224 6876
rect 11510 6872 11536 6898
rect 15788 6944 15792 6961
rect 15792 6944 15809 6961
rect 15809 6944 15814 6961
rect 15788 6940 15814 6944
rect 16294 6961 16320 6966
rect 16294 6944 16298 6961
rect 16298 6944 16315 6961
rect 16315 6944 16320 6961
rect 16294 6940 16320 6944
rect 17858 6940 17884 6966
rect 18410 6974 18436 7000
rect 20158 6974 20184 7000
rect 21308 6995 21334 7000
rect 18088 6961 18114 6966
rect 18088 6944 18092 6961
rect 18092 6944 18109 6961
rect 18109 6944 18114 6961
rect 18088 6940 18114 6944
rect 18318 6961 18344 6966
rect 18318 6944 18322 6961
rect 18322 6944 18339 6961
rect 18339 6944 18344 6961
rect 18318 6940 18344 6944
rect 19606 6940 19632 6966
rect 19882 6940 19908 6966
rect 14408 6872 14434 6898
rect 15742 6927 15768 6932
rect 15742 6910 15746 6927
rect 15746 6910 15763 6927
rect 15763 6910 15768 6927
rect 15742 6906 15768 6910
rect 16570 6906 16596 6932
rect 18870 6906 18896 6932
rect 19376 6906 19402 6932
rect 19974 6906 20000 6932
rect 20342 6961 20368 6966
rect 20342 6944 20346 6961
rect 20346 6944 20363 6961
rect 20363 6944 20368 6961
rect 20342 6940 20368 6944
rect 21078 6961 21104 6966
rect 21078 6944 21082 6961
rect 21082 6944 21099 6961
rect 21099 6944 21104 6961
rect 21078 6940 21104 6944
rect 21308 6978 21310 6995
rect 21310 6978 21334 6995
rect 21308 6974 21334 6978
rect 23516 6995 23542 7000
rect 23516 6978 23518 6995
rect 23518 6978 23542 6995
rect 23516 6974 23542 6978
rect 25954 6974 25980 7000
rect 29128 6995 29154 7000
rect 29128 6978 29132 6995
rect 29132 6978 29149 6995
rect 29149 6978 29154 6995
rect 29128 6974 29154 6978
rect 21354 6940 21380 6966
rect 22596 6961 22622 6966
rect 22596 6944 22600 6961
rect 22600 6944 22617 6961
rect 22617 6944 22622 6961
rect 22596 6940 22622 6944
rect 22642 6961 22668 6966
rect 22642 6944 22657 6961
rect 22657 6944 22668 6961
rect 22642 6940 22668 6944
rect 22734 6961 22760 6966
rect 22734 6944 22758 6961
rect 22758 6944 22760 6961
rect 22734 6940 22760 6944
rect 22918 6961 22944 6966
rect 22918 6944 22929 6961
rect 22929 6944 22944 6961
rect 22918 6940 22944 6944
rect 23240 6940 23266 6966
rect 23562 6940 23588 6966
rect 24758 6961 24784 6966
rect 24758 6944 24762 6961
rect 24762 6944 24779 6961
rect 24779 6944 24784 6961
rect 24758 6940 24784 6944
rect 24850 6961 24876 6966
rect 24850 6944 24854 6961
rect 24854 6944 24871 6961
rect 24871 6944 24876 6961
rect 24850 6940 24876 6944
rect 24896 6961 24922 6966
rect 24896 6944 24900 6961
rect 24900 6944 24917 6961
rect 24917 6944 24922 6961
rect 24896 6940 24922 6944
rect 26092 6940 26118 6966
rect 29036 6961 29062 6966
rect 29036 6944 29040 6961
rect 29040 6944 29057 6961
rect 29057 6944 29062 6961
rect 29036 6940 29062 6944
rect 29174 6961 29200 6966
rect 29174 6944 29178 6961
rect 29178 6944 29195 6961
rect 29195 6944 29200 6961
rect 29174 6940 29200 6944
rect 29358 6940 29384 6966
rect 17398 6872 17424 6898
rect 22090 6872 22116 6898
rect 22780 6872 22806 6898
rect 6220 6859 6246 6864
rect 6220 6842 6224 6859
rect 6224 6842 6241 6859
rect 6241 6842 6246 6859
rect 6220 6838 6246 6842
rect 6772 6838 6798 6864
rect 13764 6838 13790 6864
rect 24114 6838 24140 6864
rect 25678 6927 25704 6932
rect 25678 6910 25682 6927
rect 25682 6910 25699 6927
rect 25699 6910 25704 6927
rect 25678 6906 25704 6910
rect 24712 6872 24738 6898
rect 26736 6872 26762 6898
rect 29312 6893 29338 6898
rect 29312 6876 29316 6893
rect 29316 6876 29333 6893
rect 29333 6876 29338 6893
rect 29312 6872 29338 6876
rect 24574 6838 24600 6864
rect 14408 6757 14434 6762
rect 14408 6740 14412 6757
rect 14412 6740 14429 6757
rect 14429 6740 14434 6757
rect 14408 6736 14434 6740
rect 22642 6736 22668 6762
rect 24850 6736 24876 6762
rect 29036 6736 29062 6762
rect 6082 6702 6108 6728
rect 6220 6668 6246 6694
rect 10820 6689 10846 6694
rect 10820 6672 10824 6689
rect 10824 6672 10841 6689
rect 10841 6672 10846 6689
rect 10820 6668 10846 6672
rect 11142 6668 11168 6694
rect 20250 6668 20276 6694
rect 23240 6668 23266 6694
rect 23976 6689 24002 6694
rect 23976 6672 23980 6689
rect 23980 6672 23997 6689
rect 23997 6672 24002 6689
rect 23976 6668 24002 6672
rect 27978 6689 28004 6694
rect 27978 6672 27982 6689
rect 27982 6672 27999 6689
rect 27999 6672 28004 6689
rect 27978 6668 28004 6672
rect 6220 6600 6246 6626
rect 7784 6634 7810 6660
rect 13626 6634 13652 6660
rect 13764 6634 13790 6660
rect 17858 6655 17884 6660
rect 17858 6638 17862 6655
rect 17862 6638 17879 6655
rect 17879 6638 17884 6655
rect 17858 6634 17884 6638
rect 6910 6600 6936 6626
rect 11004 6600 11030 6626
rect 11832 6621 11858 6626
rect 11832 6604 11836 6621
rect 11836 6604 11853 6621
rect 11853 6604 11858 6621
rect 11832 6600 11858 6604
rect 16110 6600 16136 6626
rect 18088 6634 18114 6660
rect 18962 6655 18988 6660
rect 18962 6638 18966 6655
rect 18966 6638 18983 6655
rect 18983 6638 18988 6655
rect 18962 6634 18988 6638
rect 19146 6655 19172 6660
rect 19146 6638 19150 6655
rect 19150 6638 19167 6655
rect 19167 6638 19172 6655
rect 19146 6634 19172 6638
rect 19330 6634 19356 6660
rect 21078 6634 21104 6660
rect 21262 6634 21288 6660
rect 21354 6655 21380 6660
rect 21354 6638 21375 6655
rect 21375 6638 21380 6655
rect 21354 6634 21380 6638
rect 24114 6655 24140 6660
rect 24114 6638 24135 6655
rect 24135 6638 24140 6655
rect 24114 6634 24140 6638
rect 28392 6634 28418 6660
rect 21124 6600 21150 6626
rect 21446 6621 21472 6626
rect 21446 6604 21448 6621
rect 21448 6604 21472 6621
rect 21446 6600 21472 6604
rect 24206 6621 24232 6626
rect 24206 6604 24208 6621
rect 24208 6604 24232 6621
rect 24206 6600 24232 6604
rect 28208 6621 28234 6626
rect 28208 6604 28210 6621
rect 28210 6604 28234 6621
rect 28208 6600 28234 6604
rect 5990 6587 6016 6592
rect 5990 6570 5997 6587
rect 5997 6570 6014 6587
rect 6014 6570 6016 6587
rect 5990 6566 6016 6570
rect 6128 6566 6154 6592
rect 6726 6566 6752 6592
rect 18134 6566 18160 6592
rect 6128 6485 6154 6490
rect 6128 6468 6132 6485
rect 6132 6468 6149 6485
rect 6149 6468 6154 6485
rect 6128 6464 6154 6468
rect 6220 6430 6246 6456
rect 6496 6430 6522 6456
rect 6174 6396 6200 6422
rect 6082 6362 6108 6388
rect 5944 6328 5970 6354
rect 6726 6451 6752 6456
rect 6726 6434 6730 6451
rect 6730 6434 6747 6451
rect 6747 6434 6752 6451
rect 6726 6430 6752 6434
rect 22734 6464 22760 6490
rect 24344 6464 24370 6490
rect 7600 6430 7626 6456
rect 15926 6430 15952 6456
rect 16018 6430 16044 6456
rect 15972 6417 15998 6422
rect 15972 6400 15976 6417
rect 15976 6400 15993 6417
rect 15993 6400 15998 6417
rect 15972 6396 15998 6400
rect 16110 6417 16136 6422
rect 16110 6400 16114 6417
rect 16114 6400 16131 6417
rect 16131 6400 16136 6417
rect 16110 6396 16136 6400
rect 17858 6430 17884 6456
rect 6588 6383 6614 6388
rect 6588 6366 6592 6383
rect 6592 6366 6609 6383
rect 6609 6366 6614 6383
rect 6588 6362 6614 6366
rect 7600 6383 7626 6388
rect 7600 6366 7604 6383
rect 7604 6366 7621 6383
rect 7621 6366 7626 6383
rect 7600 6362 7626 6366
rect 16294 6362 16320 6388
rect 17122 6417 17148 6422
rect 17122 6400 17126 6417
rect 17126 6400 17143 6417
rect 17143 6400 17148 6417
rect 17122 6396 17148 6400
rect 17030 6362 17056 6388
rect 18134 6417 18160 6422
rect 18134 6400 18138 6417
rect 18138 6400 18155 6417
rect 18155 6400 18160 6417
rect 18134 6396 18160 6400
rect 19146 6430 19172 6456
rect 18410 6417 18436 6422
rect 18410 6400 18414 6417
rect 18414 6400 18431 6417
rect 18431 6400 18436 6417
rect 18410 6396 18436 6400
rect 19330 6430 19356 6456
rect 19376 6451 19402 6456
rect 19376 6434 19380 6451
rect 19380 6434 19397 6451
rect 19397 6434 19402 6451
rect 19376 6430 19402 6434
rect 18686 6362 18712 6388
rect 20112 6396 20138 6422
rect 20204 6417 20230 6422
rect 20204 6400 20208 6417
rect 20208 6400 20225 6417
rect 20225 6400 20230 6417
rect 20204 6396 20230 6400
rect 20572 6451 20598 6456
rect 20572 6434 20576 6451
rect 20576 6434 20593 6451
rect 20593 6434 20598 6451
rect 20572 6430 20598 6434
rect 21308 6451 21334 6456
rect 21308 6434 21310 6451
rect 21310 6434 21334 6451
rect 21308 6430 21334 6434
rect 23378 6451 23404 6456
rect 23378 6434 23380 6451
rect 23380 6434 23404 6451
rect 23378 6430 23404 6434
rect 24574 6451 24600 6456
rect 24574 6434 24578 6451
rect 24578 6434 24595 6451
rect 24595 6434 24600 6451
rect 24574 6430 24600 6434
rect 24758 6464 24784 6490
rect 25448 6430 25474 6456
rect 28484 6430 28510 6456
rect 21078 6417 21104 6422
rect 21078 6400 21082 6417
rect 21082 6400 21099 6417
rect 21099 6400 21104 6417
rect 21078 6396 21104 6400
rect 21354 6396 21380 6422
rect 23194 6396 23220 6422
rect 23562 6396 23588 6422
rect 5990 6294 6016 6320
rect 6266 6315 6292 6320
rect 6266 6298 6270 6315
rect 6270 6298 6287 6315
rect 6287 6298 6292 6315
rect 6266 6294 6292 6298
rect 16524 6315 16550 6320
rect 16524 6298 16528 6315
rect 16528 6298 16545 6315
rect 16545 6298 16550 6315
rect 16524 6294 16550 6298
rect 22964 6294 22990 6320
rect 27978 6396 28004 6422
rect 28208 6417 28234 6422
rect 28208 6400 28212 6417
rect 28212 6400 28229 6417
rect 28229 6400 28234 6417
rect 28208 6396 28234 6400
rect 28346 6417 28372 6422
rect 28346 6400 28367 6417
rect 28367 6400 28372 6417
rect 28346 6396 28372 6400
rect 29174 6362 29200 6388
rect 5530 6192 5556 6218
rect 6588 6192 6614 6218
rect 6910 6192 6936 6218
rect 6128 6158 6154 6184
rect 6266 6124 6292 6150
rect 5944 6056 5970 6082
rect 6496 6077 6522 6082
rect 6496 6060 6500 6077
rect 6500 6060 6517 6077
rect 6517 6060 6522 6077
rect 6496 6056 6522 6060
rect 6772 6158 6798 6184
rect 7646 6158 7672 6184
rect 7600 6124 7626 6150
rect 8014 6124 8040 6150
rect 21308 6124 21334 6150
rect 7784 6111 7810 6116
rect 7784 6094 7788 6111
rect 7788 6094 7805 6111
rect 7805 6094 7810 6111
rect 7784 6090 7810 6094
rect 11050 6090 11076 6116
rect 19882 6111 19908 6116
rect 19882 6094 19886 6111
rect 19886 6094 19903 6111
rect 19903 6094 19908 6111
rect 19882 6090 19908 6094
rect 19974 6090 20000 6116
rect 20158 6090 20184 6116
rect 7508 6043 7534 6048
rect 7508 6026 7512 6043
rect 7512 6026 7529 6043
rect 7529 6026 7534 6043
rect 7508 6022 7534 6026
rect 7646 6056 7672 6082
rect 9256 6022 9282 6048
rect 11556 6022 11582 6048
rect 7508 5920 7534 5946
rect 11096 5920 11122 5946
rect 18548 5920 18574 5946
rect 29680 5920 29706 5946
rect 7830 5886 7856 5912
rect 8244 5886 8270 5912
rect 9256 5886 9282 5912
rect 7738 5852 7764 5878
rect 9302 5873 9328 5878
rect 9302 5856 9306 5873
rect 9306 5856 9323 5873
rect 9323 5856 9328 5873
rect 9302 5852 9328 5856
rect 9486 5907 9512 5912
rect 9486 5890 9490 5907
rect 9490 5890 9507 5907
rect 9507 5890 9512 5907
rect 9486 5886 9512 5890
rect 10452 5886 10478 5912
rect 9440 5873 9466 5878
rect 9440 5856 9444 5873
rect 9444 5856 9461 5873
rect 9461 5856 9466 5873
rect 9440 5852 9466 5856
rect 9532 5873 9558 5878
rect 9532 5856 9539 5873
rect 9539 5856 9556 5873
rect 9556 5856 9558 5873
rect 9532 5852 9558 5856
rect 8106 5839 8132 5844
rect 8106 5822 8110 5839
rect 8110 5822 8127 5839
rect 8127 5822 8132 5839
rect 8106 5818 8132 5822
rect 10130 5873 10156 5878
rect 10130 5856 10134 5873
rect 10134 5856 10151 5873
rect 10151 5856 10156 5873
rect 10130 5852 10156 5856
rect 10176 5873 10202 5878
rect 10176 5856 10180 5873
rect 10180 5856 10197 5873
rect 10197 5856 10202 5873
rect 10176 5852 10202 5856
rect 11004 5818 11030 5844
rect 11556 5873 11582 5878
rect 11556 5856 11560 5873
rect 11560 5856 11577 5873
rect 11577 5856 11582 5873
rect 11556 5852 11582 5856
rect 11832 5886 11858 5912
rect 18088 5886 18114 5912
rect 17030 5852 17056 5878
rect 17122 5873 17148 5878
rect 17122 5856 17126 5873
rect 17126 5856 17143 5873
rect 17143 5856 17148 5873
rect 17122 5852 17148 5856
rect 17214 5852 17240 5878
rect 18272 5852 18298 5878
rect 18502 5852 18528 5878
rect 19100 5886 19126 5912
rect 19330 5852 19356 5878
rect 19836 5873 19862 5878
rect 19836 5856 19840 5873
rect 19840 5856 19857 5873
rect 19857 5856 19862 5873
rect 19836 5852 19862 5856
rect 20710 5886 20736 5912
rect 26230 5886 26256 5912
rect 28576 5886 28602 5912
rect 24206 5852 24232 5878
rect 28346 5852 28372 5878
rect 20112 5839 20138 5844
rect 20112 5822 20116 5839
rect 20116 5822 20133 5839
rect 20133 5822 20138 5839
rect 20112 5818 20138 5822
rect 7876 5750 7902 5776
rect 9026 5750 9052 5776
rect 11648 5771 11674 5776
rect 11648 5754 11652 5771
rect 11652 5754 11669 5771
rect 11669 5754 11674 5771
rect 11648 5750 11674 5754
rect 15926 5750 15952 5776
rect 28208 5784 28234 5810
rect 27288 5750 27314 5776
rect 10130 5648 10156 5674
rect 7876 5601 7902 5606
rect 7876 5584 7880 5601
rect 7880 5584 7897 5601
rect 7897 5584 7902 5601
rect 7876 5580 7902 5584
rect 7830 5567 7856 5572
rect 7830 5550 7834 5567
rect 7834 5550 7851 5567
rect 7851 5550 7856 5567
rect 7830 5546 7856 5550
rect 7922 5567 7948 5572
rect 7922 5550 7926 5567
rect 7926 5550 7943 5567
rect 7943 5550 7948 5567
rect 7922 5546 7948 5550
rect 8014 5567 8040 5572
rect 8014 5550 8018 5567
rect 8018 5550 8035 5567
rect 8035 5550 8040 5567
rect 8014 5546 8040 5550
rect 7738 5533 7764 5538
rect 7738 5516 7742 5533
rect 7742 5516 7759 5533
rect 7759 5516 7764 5533
rect 8612 5567 8638 5572
rect 8612 5550 8616 5567
rect 8616 5550 8633 5567
rect 8633 5550 8638 5567
rect 8612 5546 8638 5550
rect 8980 5546 9006 5572
rect 9026 5567 9052 5572
rect 9026 5550 9030 5567
rect 9030 5550 9047 5567
rect 9047 5550 9052 5567
rect 9026 5546 9052 5550
rect 16570 5614 16596 5640
rect 9486 5580 9512 5606
rect 11648 5580 11674 5606
rect 10222 5567 10248 5572
rect 10222 5550 10226 5567
rect 10226 5550 10243 5567
rect 10243 5550 10248 5567
rect 10222 5546 10248 5550
rect 16064 5580 16090 5606
rect 16524 5580 16550 5606
rect 17030 5580 17056 5606
rect 18686 5669 18712 5674
rect 18686 5652 18690 5669
rect 18690 5652 18707 5669
rect 18707 5652 18712 5669
rect 18686 5648 18712 5652
rect 19836 5669 19862 5674
rect 19836 5652 19840 5669
rect 19840 5652 19857 5669
rect 19857 5652 19862 5669
rect 19836 5648 19862 5652
rect 18502 5567 18528 5572
rect 7738 5512 7764 5516
rect 9440 5512 9466 5538
rect 15236 5512 15262 5538
rect 17122 5512 17148 5538
rect 18502 5550 18506 5567
rect 18506 5550 18523 5567
rect 18523 5550 18528 5567
rect 18502 5546 18528 5550
rect 18548 5567 18574 5572
rect 18548 5550 18552 5567
rect 18552 5550 18569 5567
rect 18569 5550 18574 5567
rect 18548 5546 18574 5550
rect 17398 5533 17424 5538
rect 17398 5516 17415 5533
rect 17415 5516 17424 5533
rect 17398 5512 17424 5516
rect 18272 5512 18298 5538
rect 19606 5546 19632 5572
rect 19974 5580 20000 5606
rect 19882 5546 19908 5572
rect 22136 5567 22162 5572
rect 22136 5550 22140 5567
rect 22140 5550 22157 5567
rect 22157 5550 22162 5567
rect 22136 5546 22162 5550
rect 22274 5614 22300 5640
rect 25402 5614 25428 5640
rect 27012 5580 27038 5606
rect 22274 5567 22300 5572
rect 22274 5550 22298 5567
rect 22298 5550 22300 5567
rect 22274 5546 22300 5550
rect 21952 5512 21978 5538
rect 22688 5546 22714 5572
rect 25356 5546 25382 5572
rect 25678 5512 25704 5538
rect 26828 5512 26854 5538
rect 27104 5546 27130 5572
rect 27288 5567 27314 5572
rect 27288 5550 27292 5567
rect 27292 5550 27309 5567
rect 27309 5550 27314 5567
rect 27288 5546 27314 5550
rect 10176 5478 10202 5504
rect 15696 5499 15722 5504
rect 15696 5482 15700 5499
rect 15700 5482 15717 5499
rect 15717 5482 15722 5499
rect 15696 5478 15722 5482
rect 16984 5499 17010 5504
rect 16984 5482 16988 5499
rect 16988 5482 17005 5499
rect 17005 5482 17010 5499
rect 16984 5478 17010 5482
rect 22320 5478 22346 5504
rect 22412 5478 22438 5504
rect 8014 5376 8040 5402
rect 9532 5376 9558 5402
rect 11004 5376 11030 5402
rect 15972 5397 15998 5402
rect 15972 5380 15976 5397
rect 15976 5380 15993 5397
rect 15993 5380 15998 5397
rect 15972 5376 15998 5380
rect 16064 5397 16090 5402
rect 16064 5380 16068 5397
rect 16068 5380 16085 5397
rect 16085 5380 16090 5397
rect 16064 5376 16090 5380
rect 17398 5397 17424 5402
rect 17398 5380 17402 5397
rect 17402 5380 17419 5397
rect 17419 5380 17424 5397
rect 17398 5376 17424 5380
rect 22274 5376 22300 5402
rect 25356 5397 25382 5402
rect 25356 5380 25360 5397
rect 25360 5380 25377 5397
rect 25377 5380 25382 5397
rect 25356 5376 25382 5380
rect 25448 5376 25474 5402
rect 7738 5342 7764 5368
rect 7922 5308 7948 5334
rect 8290 5329 8316 5334
rect 8290 5312 8294 5329
rect 8294 5312 8311 5329
rect 8311 5312 8316 5329
rect 8290 5308 8316 5312
rect 8244 5274 8270 5300
rect 9440 5308 9466 5334
rect 15696 5342 15722 5368
rect 13626 5308 13652 5334
rect 17122 5342 17148 5368
rect 15926 5329 15952 5334
rect 15926 5312 15930 5329
rect 15930 5312 15947 5329
rect 15947 5312 15952 5329
rect 15926 5308 15952 5312
rect 16110 5329 16136 5334
rect 16110 5312 16114 5329
rect 16114 5312 16131 5329
rect 16131 5312 16136 5329
rect 16110 5308 16136 5312
rect 16984 5308 17010 5334
rect 20112 5342 20138 5368
rect 20848 5342 20874 5368
rect 21308 5363 21334 5368
rect 21308 5346 21310 5363
rect 21310 5346 21334 5363
rect 21308 5342 21334 5346
rect 23378 5342 23404 5368
rect 18272 5308 18298 5334
rect 18962 5308 18988 5334
rect 20158 5329 20184 5334
rect 20158 5312 20162 5329
rect 20162 5312 20179 5329
rect 20179 5312 20184 5329
rect 20158 5308 20184 5312
rect 21078 5329 21104 5334
rect 21078 5312 21082 5329
rect 21082 5312 21099 5329
rect 21099 5312 21104 5329
rect 21078 5308 21104 5312
rect 21354 5308 21380 5334
rect 23838 5308 23864 5334
rect 24206 5308 24232 5334
rect 25356 5329 25382 5334
rect 25356 5312 25360 5329
rect 25360 5312 25377 5329
rect 25377 5312 25382 5329
rect 25356 5308 25382 5312
rect 25402 5329 25428 5334
rect 25402 5312 25417 5329
rect 25417 5312 25428 5329
rect 25402 5308 25428 5312
rect 25678 5329 25704 5334
rect 25678 5312 25689 5329
rect 25689 5312 25704 5329
rect 16018 5295 16044 5300
rect 16018 5278 16022 5295
rect 16022 5278 16039 5295
rect 16039 5278 16044 5295
rect 16018 5274 16044 5278
rect 10222 5240 10248 5266
rect 18318 5295 18344 5300
rect 8290 5206 8316 5232
rect 8612 5206 8638 5232
rect 16018 5206 16044 5232
rect 18318 5278 18322 5295
rect 18322 5278 18339 5295
rect 18339 5278 18344 5295
rect 18318 5274 18344 5278
rect 17030 5240 17056 5266
rect 25678 5308 25704 5312
rect 25632 5240 25658 5266
rect 18640 5206 18666 5232
rect 20848 5206 20874 5232
rect 23378 5206 23404 5232
rect 8290 5104 8316 5130
rect 22136 5104 22162 5130
rect 25356 5104 25382 5130
rect 18272 5036 18298 5062
rect 7830 5002 7856 5028
rect 8244 5002 8270 5028
rect 18962 5036 18988 5062
rect 21078 5036 21104 5062
rect 23838 5036 23864 5062
rect 18640 5023 18666 5028
rect 18640 5006 18644 5023
rect 18644 5006 18661 5023
rect 18661 5006 18666 5023
rect 18640 5002 18666 5006
rect 19606 5023 19632 5028
rect 19606 5006 19610 5023
rect 19610 5006 19627 5023
rect 19627 5006 19632 5023
rect 19606 5002 19632 5006
rect 19882 5002 19908 5028
rect 21354 5023 21380 5028
rect 21354 5006 21375 5023
rect 21375 5006 21380 5023
rect 21354 5002 21380 5006
rect 24252 5002 24278 5028
rect 21446 4989 21472 4994
rect 21446 4972 21448 4989
rect 21448 4972 21472 4989
rect 21446 4968 21472 4972
rect 24206 4989 24232 4994
rect 24206 4972 24208 4989
rect 24208 4972 24232 4989
rect 24206 4968 24232 4972
rect 18456 4934 18482 4960
rect 18594 4955 18620 4960
rect 18594 4938 18598 4955
rect 18598 4938 18615 4955
rect 18615 4938 18620 4955
rect 18594 4934 18620 4938
rect 15972 4832 15998 4858
rect 15926 4798 15952 4824
rect 18318 4832 18344 4858
rect 17260 4798 17286 4824
rect 18594 4798 18620 4824
rect 17030 4764 17056 4790
rect 17214 4785 17240 4790
rect 17214 4768 17218 4785
rect 17218 4768 17235 4785
rect 17235 4768 17240 4785
rect 17214 4764 17240 4768
rect 18456 4764 18482 4790
rect 19606 4798 19632 4824
rect 17122 4730 17148 4756
rect 19882 4764 19908 4790
rect 21124 4798 21150 4824
rect 22412 4798 22438 4824
rect 21078 4785 21104 4790
rect 21078 4768 21082 4785
rect 21082 4768 21099 4785
rect 21099 4768 21104 4785
rect 21078 4764 21104 4768
rect 21354 4764 21380 4790
rect 17076 4683 17102 4688
rect 17076 4666 17080 4683
rect 17080 4666 17097 4683
rect 17097 4666 17102 4683
rect 17076 4662 17102 4666
rect 17122 4560 17148 4586
rect 17260 4581 17286 4586
rect 17260 4564 17264 4581
rect 17264 4564 17281 4581
rect 17281 4564 17286 4581
rect 17260 4560 17286 4564
rect 19606 4560 19632 4586
rect 25632 4560 25658 4586
rect 23838 4492 23864 4518
rect 17076 4458 17102 4484
rect 24206 4479 24232 4484
rect 24206 4462 24227 4479
rect 24227 4462 24232 4479
rect 24206 4458 24232 4462
rect 21124 4424 21150 4450
rect 25954 4458 25980 4484
rect 18640 3969 18666 3974
rect 18640 3952 18644 3969
rect 18644 3952 18661 3969
rect 18661 3952 18666 3969
rect 18640 3948 18666 3952
rect 19192 3948 19218 3974
rect 18778 3935 18804 3940
rect 18778 3918 18782 3935
rect 18782 3918 18799 3935
rect 18799 3918 18804 3935
rect 18778 3914 18804 3918
rect 20388 3914 20414 3940
rect 16294 650 16320 676
rect 16708 650 16734 676
<< metal2 >>
rect 4702 28964 4728 28967
rect 4702 28935 4728 28938
rect 4708 28695 4722 28935
rect 4932 28930 4958 28933
rect 4932 28901 4958 28904
rect 4702 28692 4728 28695
rect 4702 28663 4728 28666
rect 4518 27604 4544 27607
rect 4518 27575 4544 27578
rect 4524 27335 4538 27575
rect 4708 27335 4722 28663
rect 4938 28253 4952 28901
rect 5536 28797 5550 33000
rect 5576 28930 5602 28933
rect 5576 28901 5602 28904
rect 5530 28794 5556 28797
rect 5530 28765 5556 28768
rect 5162 28692 5188 28695
rect 5162 28663 5188 28666
rect 5168 28525 5182 28663
rect 5162 28522 5188 28525
rect 5162 28493 5188 28496
rect 5484 28454 5510 28457
rect 5484 28425 5510 28428
rect 4932 28250 4958 28253
rect 4932 28221 4958 28224
rect 5490 28151 5504 28425
rect 5536 28423 5550 28765
rect 5582 28729 5596 28901
rect 5628 28899 5642 33000
rect 14230 32968 14336 32982
rect 10268 29576 10294 29579
rect 10268 29547 10294 29550
rect 8704 29474 8730 29477
rect 8704 29445 8730 29448
rect 7048 29304 7074 29307
rect 7048 29275 7074 29278
rect 6956 29270 6982 29273
rect 6956 29241 6982 29244
rect 6726 29236 6752 29239
rect 6726 29207 6752 29210
rect 5622 28896 5648 28899
rect 5622 28867 5648 28870
rect 5576 28726 5602 28729
rect 5576 28697 5602 28700
rect 5530 28420 5556 28423
rect 5530 28391 5556 28394
rect 5530 28352 5556 28355
rect 5530 28323 5556 28326
rect 5484 28148 5510 28151
rect 5484 28119 5510 28122
rect 4794 27672 4820 27675
rect 4794 27643 4820 27646
rect 4518 27332 4544 27335
rect 4518 27303 4544 27306
rect 4702 27332 4728 27335
rect 4702 27303 4728 27306
rect 4524 27063 4538 27303
rect 4800 27097 4814 27643
rect 5070 27638 5096 27641
rect 5070 27609 5096 27612
rect 4656 27094 4682 27097
rect 4656 27065 4682 27068
rect 4794 27094 4820 27097
rect 4794 27065 4820 27068
rect 4518 27060 4544 27063
rect 4518 27031 4544 27034
rect 4472 26040 4498 26043
rect 4472 26011 4498 26014
rect 3276 25496 3302 25499
rect 3276 25467 3302 25470
rect 3282 25159 3296 25467
rect 3414 25462 3440 25465
rect 3414 25433 3440 25436
rect 3644 25462 3670 25465
rect 3644 25433 3670 25436
rect 3420 25261 3434 25433
rect 3414 25258 3440 25261
rect 3414 25229 3440 25232
rect 3276 25156 3302 25159
rect 3276 25127 3302 25130
rect 3282 24377 3296 25127
rect 3276 24374 3302 24377
rect 3276 24345 3302 24348
rect 3420 24343 3434 25229
rect 3506 24374 3532 24377
rect 3506 24345 3532 24348
rect 3414 24340 3440 24343
rect 3414 24311 3440 24314
rect 3420 24173 3434 24311
rect 3414 24170 3440 24173
rect 3414 24141 3440 24144
rect 3367 24052 3395 24056
rect 3184 24034 3210 24037
rect 3367 24019 3368 24024
rect 3184 24005 3210 24008
rect 3394 24019 3395 24024
rect 3368 24005 3394 24008
rect 3138 22436 3164 22439
rect 3138 22407 3164 22410
rect 3144 22167 3158 22407
rect 3190 22405 3204 24005
rect 3420 23799 3434 24141
rect 3512 24113 3526 24345
rect 3466 24099 3526 24113
rect 3466 24071 3480 24099
rect 3460 24068 3486 24071
rect 3460 24039 3486 24042
rect 3466 23867 3480 24039
rect 3460 23864 3486 23867
rect 3460 23835 3486 23838
rect 3414 23796 3440 23799
rect 3414 23767 3440 23770
rect 3420 23527 3434 23767
rect 3414 23524 3440 23527
rect 3414 23495 3440 23498
rect 3466 23493 3480 23835
rect 3650 23731 3664 25433
rect 4478 25397 4492 26011
rect 4524 25907 4538 27031
rect 4518 25904 4544 25907
rect 4518 25875 4544 25878
rect 4472 25394 4498 25397
rect 4472 25365 4498 25368
rect 3736 25156 3762 25159
rect 3736 25127 3762 25130
rect 3690 23864 3716 23867
rect 3690 23835 3716 23838
rect 3644 23728 3670 23731
rect 3644 23699 3670 23702
rect 3460 23490 3486 23493
rect 3460 23461 3486 23464
rect 3552 22742 3578 22745
rect 3552 22713 3578 22716
rect 3414 22708 3440 22711
rect 3414 22679 3440 22682
rect 3184 22402 3210 22405
rect 3184 22373 3210 22376
rect 3190 22345 3204 22373
rect 3190 22331 3388 22345
rect 3138 22164 3164 22167
rect 3138 22135 3164 22138
rect 3184 21144 3210 21147
rect 3184 21115 3210 21118
rect 3190 20773 3204 21115
rect 3184 20770 3210 20773
rect 3184 20741 3210 20744
rect 3138 19172 3164 19175
rect 3138 19143 3164 19146
rect 3144 18937 3158 19143
rect 3374 19141 3388 22331
rect 3420 22167 3434 22679
rect 3558 22439 3572 22713
rect 3552 22436 3578 22439
rect 3552 22407 3578 22410
rect 3558 22201 3572 22407
rect 3552 22198 3578 22201
rect 3552 22169 3578 22172
rect 3414 22164 3440 22167
rect 3414 22135 3440 22138
rect 3420 21623 3434 22135
rect 3460 21688 3486 21691
rect 3460 21659 3486 21662
rect 3414 21620 3440 21623
rect 3414 21591 3440 21594
rect 3420 21113 3434 21591
rect 3414 21110 3440 21113
rect 3414 21081 3440 21084
rect 3414 20906 3440 20909
rect 3414 20877 3440 20880
rect 3420 20773 3434 20877
rect 3414 20770 3440 20773
rect 3414 20741 3440 20744
rect 3368 19138 3394 19141
rect 3368 19109 3394 19112
rect 3374 19081 3388 19109
rect 3328 19067 3388 19081
rect 3138 18934 3164 18937
rect 3138 18905 3164 18908
rect 3144 18393 3158 18905
rect 3138 18390 3164 18393
rect 3138 18361 3164 18364
rect 3144 18087 3158 18361
rect 3138 18084 3164 18087
rect 3138 18055 3164 18058
rect 3144 17577 3158 18055
rect 3138 17574 3164 17577
rect 3138 17545 3164 17548
rect 3144 17271 3158 17545
rect 3184 17540 3210 17543
rect 3184 17511 3210 17514
rect 3138 17268 3164 17271
rect 3138 17239 3164 17242
rect 3144 16236 3158 17239
rect 3137 16232 3165 16236
rect 3137 16199 3138 16204
rect 3164 16199 3165 16204
rect 3138 16185 3164 16188
rect 3144 15945 3158 16185
rect 3138 15942 3164 15945
rect 3138 15913 3164 15916
rect 3144 15639 3158 15913
rect 3138 15636 3164 15639
rect 3138 15607 3164 15610
rect 3190 14823 3204 17511
rect 3328 15877 3342 19067
rect 3420 17509 3434 20741
rect 3466 20707 3480 21659
rect 3558 21657 3572 22169
rect 3650 21691 3664 23699
rect 3696 22745 3710 23835
rect 3690 22742 3716 22745
rect 3690 22713 3716 22716
rect 3644 21688 3670 21691
rect 3644 21659 3670 21662
rect 3552 21654 3578 21657
rect 3552 21625 3578 21628
rect 3558 21181 3572 21625
rect 3696 21453 3710 22713
rect 3690 21450 3716 21453
rect 3690 21421 3716 21424
rect 3552 21178 3578 21181
rect 3552 21149 3578 21152
rect 3552 21110 3578 21113
rect 3552 21081 3578 21084
rect 3558 20807 3572 21081
rect 3552 20804 3578 20807
rect 3552 20775 3578 20778
rect 3466 20693 3526 20707
rect 3512 18401 3526 20693
rect 3558 20569 3572 20775
rect 3552 20566 3578 20569
rect 3552 20537 3578 20540
rect 3558 20263 3572 20537
rect 3552 20260 3578 20263
rect 3552 20231 3578 20234
rect 3558 19481 3572 20231
rect 3552 19478 3578 19481
rect 3552 19449 3578 19452
rect 3598 19478 3624 19481
rect 3598 19449 3624 19452
rect 3552 19172 3578 19175
rect 3604 19149 3618 19449
rect 3578 19146 3618 19149
rect 3552 19143 3618 19146
rect 3558 19135 3618 19143
rect 3552 18934 3578 18937
rect 3604 18928 3618 19135
rect 3696 18971 3710 21421
rect 3742 21147 3756 25127
rect 3782 22198 3808 22201
rect 3782 22169 3808 22172
rect 3736 21144 3762 21147
rect 3736 21115 3762 21118
rect 3690 18968 3716 18971
rect 3690 18939 3716 18942
rect 3578 18914 3618 18928
rect 3552 18905 3578 18908
rect 3552 18424 3578 18427
rect 3512 18398 3552 18401
rect 3512 18395 3578 18398
rect 3512 18387 3572 18395
rect 3604 18393 3618 18914
rect 3598 18390 3624 18393
rect 3414 17506 3440 17509
rect 3414 17477 3440 17480
rect 3368 16214 3394 16217
rect 3394 16194 3434 16208
rect 3368 16185 3394 16188
rect 3420 15911 3434 16194
rect 3414 15908 3440 15911
rect 3414 15879 3440 15882
rect 3328 15874 3394 15877
rect 3328 15863 3368 15874
rect 3368 15845 3394 15848
rect 3420 15673 3434 15879
rect 3414 15670 3440 15673
rect 3414 15641 3440 15644
rect 3460 15636 3486 15639
rect 3460 15607 3486 15610
rect 3414 15126 3440 15129
rect 3414 15097 3440 15100
rect 3322 14922 3348 14925
rect 3322 14893 3348 14896
rect 3184 14820 3210 14823
rect 3184 14791 3210 14794
rect 3184 14752 3210 14755
rect 3184 14723 3210 14726
rect 3190 14585 3204 14723
rect 3184 14582 3210 14585
rect 3184 14553 3210 14556
rect 3190 14279 3204 14553
rect 3328 14551 3342 14893
rect 3368 14786 3394 14789
rect 3368 14757 3394 14760
rect 3322 14548 3348 14551
rect 3322 14519 3348 14522
rect 3328 14381 3342 14519
rect 3322 14378 3348 14381
rect 3322 14349 3348 14352
rect 3184 14276 3210 14279
rect 3184 14247 3210 14250
rect 3190 14075 3204 14247
rect 3184 14072 3210 14075
rect 3184 14043 3210 14046
rect 3328 14007 3342 14349
rect 3322 14004 3348 14007
rect 3322 13975 3348 13978
rect 3328 13497 3342 13975
rect 3322 13494 3348 13497
rect 3322 13465 3348 13468
rect 3328 13293 3342 13465
rect 3322 13290 3348 13293
rect 3322 13261 3348 13264
rect 3138 13222 3164 13225
rect 3138 13193 3164 13196
rect 3144 12919 3158 13193
rect 3374 13157 3388 14757
rect 3420 14585 3434 15097
rect 3466 15095 3480 15607
rect 3460 15092 3486 15095
rect 3460 15063 3486 15066
rect 3466 14925 3480 15063
rect 3460 14922 3486 14925
rect 3460 14893 3486 14896
rect 3414 14582 3440 14585
rect 3414 14553 3440 14556
rect 3460 14276 3486 14279
rect 3512 14270 3526 18387
rect 3598 18361 3624 18364
rect 3604 18189 3618 18361
rect 3598 18186 3624 18189
rect 3598 18157 3624 18160
rect 3696 16421 3710 18939
rect 3742 18087 3756 21115
rect 3788 19515 3802 22169
rect 3920 21110 3946 21113
rect 3920 21081 3946 21084
rect 3926 20739 3940 21081
rect 3920 20736 3946 20739
rect 3920 20707 3946 20710
rect 3828 20600 3854 20603
rect 3828 20571 3854 20574
rect 3782 19512 3808 19515
rect 3782 19483 3808 19486
rect 3736 18084 3762 18087
rect 3736 18055 3762 18058
rect 3690 16418 3716 16421
rect 3690 16389 3716 16392
rect 3696 15877 3710 16389
rect 3650 15863 3710 15877
rect 3742 15877 3756 18055
rect 3834 17339 3848 20571
rect 3926 20569 3940 20707
rect 4478 20569 4492 25365
rect 4662 23518 4676 27065
rect 4840 26006 4866 26009
rect 4840 25977 4866 25980
rect 4702 25904 4728 25907
rect 4702 25875 4728 25878
rect 4708 25703 4722 25875
rect 4846 25813 4860 25977
rect 4800 25799 4860 25813
rect 4800 25703 4814 25799
rect 4702 25700 4728 25703
rect 4702 25671 4728 25674
rect 4794 25700 4820 25703
rect 4794 25671 4820 25674
rect 4708 25541 4722 25671
rect 4708 25537 4860 25541
rect 4708 25533 4906 25537
rect 4708 25530 4912 25533
rect 4708 25527 4886 25530
rect 4846 25523 4886 25527
rect 4886 25501 4912 25504
rect 4794 25360 4820 25363
rect 4794 25331 4820 25334
rect 4800 25159 4814 25331
rect 4794 25156 4820 25159
rect 4794 25127 4820 25130
rect 4886 25122 4912 25125
rect 4886 25093 4912 25096
rect 4892 24668 4906 25093
rect 4885 24664 4913 24668
rect 4885 24631 4913 24636
rect 5024 24272 5050 24275
rect 5024 24243 5050 24246
rect 4932 24068 4958 24071
rect 4932 24039 4958 24042
rect 4748 24000 4774 24003
rect 4748 23971 4774 23974
rect 4754 23833 4768 23971
rect 4938 23901 4952 24039
rect 5030 23901 5044 24243
rect 5076 24139 5090 27609
rect 5254 27094 5280 27097
rect 5280 27074 5320 27088
rect 5254 27065 5280 27068
rect 5208 25700 5234 25703
rect 5208 25671 5234 25674
rect 5115 24664 5143 24668
rect 5115 24631 5143 24636
rect 5070 24136 5096 24139
rect 5070 24107 5096 24110
rect 4840 23898 4866 23901
rect 4840 23869 4866 23872
rect 4932 23898 4958 23901
rect 4932 23869 4958 23872
rect 5024 23898 5050 23901
rect 5024 23869 5050 23872
rect 4748 23830 4774 23833
rect 4748 23801 4774 23804
rect 4662 23504 4722 23518
rect 4656 22368 4682 22371
rect 4656 22339 4682 22342
rect 4662 21691 4676 22339
rect 4656 21688 4682 21691
rect 4656 21659 4682 21662
rect 4708 21589 4722 23504
rect 4846 23017 4860 23869
rect 4886 23762 4912 23765
rect 4886 23733 4912 23736
rect 4840 23014 4866 23017
rect 4840 22985 4866 22988
rect 4794 22640 4820 22643
rect 4794 22611 4820 22614
rect 4800 22439 4814 22611
rect 4846 22507 4860 22985
rect 4840 22504 4866 22507
rect 4840 22475 4866 22478
rect 4892 22473 4906 23733
rect 5070 23626 5096 23629
rect 5070 23597 5096 23600
rect 4932 22504 4958 22507
rect 4932 22475 4958 22478
rect 4886 22470 4912 22473
rect 4886 22441 4912 22444
rect 4794 22436 4820 22439
rect 4794 22407 4820 22410
rect 4748 22368 4774 22371
rect 4938 22362 4952 22475
rect 5024 22470 5050 22473
rect 5024 22441 5050 22444
rect 4978 22436 5004 22439
rect 4977 22420 4978 22424
rect 5004 22420 5005 22424
rect 4977 22387 5005 22392
rect 4938 22348 4998 22362
rect 4748 22339 4774 22342
rect 4754 22269 4768 22339
rect 4748 22266 4774 22269
rect 4748 22237 4774 22240
rect 4932 21892 4958 21895
rect 4932 21863 4958 21866
rect 4840 21654 4866 21657
rect 4840 21625 4866 21628
rect 4886 21654 4912 21657
rect 4886 21625 4912 21628
rect 4702 21586 4728 21589
rect 4702 21557 4728 21560
rect 4794 21552 4820 21555
rect 4794 21523 4820 21526
rect 4800 21317 4814 21523
rect 4656 21314 4682 21317
rect 4656 21285 4682 21288
rect 4748 21314 4774 21317
rect 4748 21285 4774 21288
rect 4794 21314 4820 21317
rect 4794 21285 4820 21288
rect 4662 20909 4676 21285
rect 4754 21147 4768 21285
rect 4748 21144 4774 21147
rect 4748 21115 4774 21118
rect 4656 20906 4682 20909
rect 4656 20877 4682 20880
rect 3920 20566 3946 20569
rect 3920 20537 3946 20540
rect 4472 20566 4498 20569
rect 4472 20537 4498 20540
rect 4702 18900 4728 18903
rect 4702 18871 4728 18874
rect 4656 18594 4682 18597
rect 4656 18565 4682 18568
rect 4662 18189 4676 18565
rect 4656 18186 4682 18189
rect 4656 18157 4682 18160
rect 4708 17645 4722 18871
rect 4702 17642 4728 17645
rect 4702 17613 4728 17616
rect 4754 17543 4768 21115
rect 4846 21045 4860 21625
rect 4892 21419 4906 21625
rect 4886 21416 4912 21419
rect 4886 21387 4912 21390
rect 4938 21385 4952 21863
rect 4932 21382 4958 21385
rect 4932 21353 4958 21356
rect 4932 21110 4958 21113
rect 4932 21081 4958 21084
rect 4840 21042 4866 21045
rect 4840 21013 4866 21016
rect 4938 20637 4952 21081
rect 4932 20634 4958 20637
rect 4932 20605 4958 20608
rect 4984 20577 4998 22348
rect 4938 20563 4998 20577
rect 4938 19481 4952 20563
rect 4978 19512 5004 19515
rect 4978 19483 5004 19486
rect 4840 19478 4866 19481
rect 4840 19449 4866 19452
rect 4932 19478 4958 19481
rect 4932 19449 4958 19452
rect 4846 19421 4860 19449
rect 4931 19428 4959 19432
rect 4846 19407 4906 19421
rect 4840 19376 4866 19379
rect 4840 19347 4866 19350
rect 4846 19005 4860 19347
rect 4892 19277 4906 19407
rect 4931 19395 4932 19400
rect 4958 19395 4959 19400
rect 4932 19381 4958 19384
rect 4886 19274 4912 19277
rect 4886 19245 4912 19248
rect 4840 19002 4866 19005
rect 4840 18973 4866 18976
rect 4840 18934 4866 18937
rect 4840 18905 4866 18908
rect 4846 18733 4860 18905
rect 4984 18835 4998 19483
rect 5030 19447 5044 22441
rect 5076 21351 5090 23597
rect 5070 21348 5096 21351
rect 5070 21319 5096 21322
rect 5024 19444 5050 19447
rect 5024 19415 5050 19418
rect 4978 18832 5004 18835
rect 4978 18803 5004 18806
rect 4840 18730 4866 18733
rect 4840 18701 4866 18704
rect 4794 18594 4820 18597
rect 4794 18565 4820 18568
rect 4800 18461 4814 18565
rect 4839 18544 4867 18548
rect 4839 18511 4867 18516
rect 4846 18461 4860 18511
rect 4794 18458 4820 18461
rect 4794 18429 4820 18432
rect 4840 18458 4866 18461
rect 4840 18429 4866 18432
rect 5030 18412 5044 19415
rect 5076 18631 5090 21319
rect 5122 21079 5136 24631
rect 5162 24612 5188 24615
rect 5214 24600 5228 25671
rect 5254 25156 5280 25159
rect 5254 25127 5280 25130
rect 5162 24583 5188 24586
rect 5207 24596 5235 24600
rect 5168 23527 5182 24583
rect 5207 24563 5235 24568
rect 5162 23524 5188 23527
rect 5162 23495 5188 23498
rect 5168 22983 5182 23495
rect 5162 22980 5188 22983
rect 5162 22951 5188 22954
rect 5161 22420 5189 22424
rect 5161 22387 5189 22392
rect 5116 21076 5142 21079
rect 5116 21047 5142 21050
rect 5070 18628 5096 18631
rect 5070 18599 5096 18602
rect 5023 18408 5051 18412
rect 5023 18375 5051 18380
rect 4748 17540 4774 17543
rect 4748 17511 4774 17514
rect 4794 17506 4820 17509
rect 4794 17477 4820 17480
rect 4800 17373 4814 17477
rect 4794 17370 4820 17373
rect 4794 17341 4820 17344
rect 3828 17336 3854 17339
rect 3828 17307 3854 17310
rect 5030 16659 5044 18375
rect 4748 16656 4774 16659
rect 4748 16627 4774 16630
rect 5024 16656 5050 16659
rect 5024 16627 5050 16630
rect 4754 16557 4768 16627
rect 4748 16554 4774 16557
rect 4748 16525 4774 16528
rect 4702 16520 4728 16523
rect 4702 16491 4728 16494
rect 4656 16452 4682 16455
rect 4656 16423 4682 16426
rect 4564 16418 4590 16421
rect 4564 16389 4590 16392
rect 4610 16418 4636 16421
rect 4610 16389 4636 16392
rect 4287 16300 4315 16304
rect 4287 16267 4288 16272
rect 4314 16267 4315 16272
rect 4288 16253 4314 16256
rect 4570 16251 4584 16389
rect 4564 16248 4590 16251
rect 4517 16232 4545 16236
rect 4472 16214 4498 16217
rect 4564 16219 4590 16222
rect 4517 16199 4518 16204
rect 4472 16185 4498 16188
rect 4544 16199 4545 16204
rect 4518 16185 4544 16188
rect 4478 16106 4492 16185
rect 4518 16112 4544 16115
rect 4478 16092 4518 16106
rect 4518 16083 4544 16086
rect 3742 15863 3802 15877
rect 3650 15698 3664 15863
rect 3690 15704 3716 15707
rect 3650 15684 3690 15698
rect 3690 15675 3716 15678
rect 3788 15163 3802 15863
rect 4616 15741 4630 16389
rect 4662 16013 4676 16423
rect 4656 16010 4682 16013
rect 4656 15981 4682 15984
rect 4610 15738 4636 15741
rect 4610 15709 4636 15712
rect 3782 15160 3808 15163
rect 3782 15131 3808 15134
rect 4708 15061 4722 16491
rect 4748 16452 4774 16455
rect 4747 16436 4748 16440
rect 4917 16452 4943 16455
rect 4774 16436 4775 16440
rect 4943 16426 4952 16446
rect 4917 16423 4952 16426
rect 4747 16403 4775 16408
rect 4938 16304 4952 16423
rect 4931 16300 4959 16304
rect 5030 16285 5044 16627
rect 4931 16267 4959 16272
rect 5024 16282 5050 16285
rect 5024 16253 5050 16256
rect 4794 16214 4820 16217
rect 4794 16185 4820 16188
rect 4800 15911 4814 16185
rect 4794 15908 4820 15911
rect 4794 15879 4820 15882
rect 5076 15129 5090 18599
rect 5122 18563 5136 21047
rect 5168 19481 5182 22387
rect 5214 22201 5228 24563
rect 5260 23731 5274 25127
rect 5254 23728 5280 23731
rect 5254 23699 5280 23702
rect 5260 23629 5274 23699
rect 5254 23626 5280 23629
rect 5254 23597 5280 23600
rect 5306 23569 5320 27074
rect 5260 23555 5320 23569
rect 5260 22949 5274 23555
rect 5346 23490 5372 23493
rect 5346 23461 5372 23464
rect 5300 22980 5326 22983
rect 5300 22951 5326 22954
rect 5254 22946 5280 22949
rect 5254 22917 5280 22920
rect 5306 22439 5320 22951
rect 5300 22436 5326 22439
rect 5300 22407 5326 22410
rect 5208 22198 5234 22201
rect 5208 22169 5234 22172
rect 5306 21997 5320 22407
rect 5352 21997 5366 23461
rect 5490 23076 5504 28119
rect 5536 27607 5550 28323
rect 5628 28253 5642 28867
rect 5990 28760 6016 28763
rect 6680 28760 6706 28763
rect 5990 28731 6016 28734
rect 6587 28744 6615 28748
rect 5622 28250 5648 28253
rect 5622 28221 5648 28224
rect 5576 28182 5602 28185
rect 5576 28153 5602 28156
rect 5530 27604 5556 27607
rect 5530 27575 5556 27578
rect 5582 27165 5596 28153
rect 5622 27298 5648 27301
rect 5622 27269 5648 27272
rect 5576 27162 5602 27165
rect 5576 27133 5602 27136
rect 5628 27131 5642 27269
rect 5622 27128 5648 27131
rect 5622 27099 5648 27102
rect 5628 26272 5642 27099
rect 5852 26448 5878 26451
rect 5852 26419 5878 26422
rect 5582 26258 5642 26272
rect 5530 26244 5556 26247
rect 5530 26215 5556 26218
rect 5536 25941 5550 26215
rect 5582 26213 5596 26258
rect 5858 26247 5872 26419
rect 5852 26244 5878 26247
rect 5852 26215 5878 26218
rect 5576 26210 5602 26213
rect 5576 26181 5602 26184
rect 5530 25938 5556 25941
rect 5530 25909 5556 25912
rect 5536 25533 5550 25909
rect 5530 25530 5556 25533
rect 5530 25501 5556 25504
rect 5536 25465 5550 25501
rect 5530 25462 5556 25465
rect 5530 25433 5556 25436
rect 5536 24615 5550 25433
rect 5806 24918 5832 24921
rect 5806 24889 5832 24892
rect 5812 24717 5826 24889
rect 5806 24714 5832 24717
rect 5806 24685 5832 24688
rect 5530 24612 5556 24615
rect 5530 24583 5556 24586
rect 5668 24612 5694 24615
rect 5668 24583 5694 24586
rect 5674 24139 5688 24583
rect 5530 24136 5556 24139
rect 5530 24107 5556 24110
rect 5668 24136 5694 24139
rect 5668 24107 5694 24110
rect 5536 23527 5550 24107
rect 5576 24000 5602 24003
rect 5576 23971 5602 23974
rect 5582 23629 5596 23971
rect 5576 23626 5602 23629
rect 5576 23597 5602 23600
rect 5530 23524 5556 23527
rect 5530 23495 5556 23498
rect 5398 23062 5504 23076
rect 5300 21994 5326 21997
rect 5300 21965 5326 21968
rect 5346 21994 5372 21997
rect 5346 21965 5372 21968
rect 5352 21937 5366 21965
rect 5214 21923 5366 21937
rect 5214 21861 5228 21923
rect 5208 21858 5234 21861
rect 5208 21829 5234 21832
rect 5346 21348 5372 21351
rect 5346 21319 5372 21322
rect 5208 21110 5234 21113
rect 5208 21081 5234 21084
rect 5162 19478 5188 19481
rect 5162 19449 5188 19452
rect 5116 18560 5142 18563
rect 5116 18531 5142 18534
rect 5214 17543 5228 21081
rect 5352 20807 5366 21319
rect 5346 20804 5372 20807
rect 5346 20775 5372 20778
rect 5352 20263 5366 20775
rect 5346 20260 5372 20263
rect 5346 20231 5372 20234
rect 5352 19753 5366 20231
rect 5346 19750 5372 19753
rect 5346 19721 5372 19724
rect 5254 18560 5280 18563
rect 5254 18531 5280 18534
rect 5208 17540 5234 17543
rect 5208 17511 5234 17514
rect 5208 15874 5234 15877
rect 5208 15845 5234 15848
rect 5214 15741 5228 15845
rect 5208 15738 5234 15741
rect 5208 15709 5234 15712
rect 5162 15160 5188 15163
rect 5162 15131 5188 15134
rect 4840 15126 4866 15129
rect 4840 15097 4866 15100
rect 4978 15126 5004 15129
rect 4978 15097 5004 15100
rect 5070 15126 5096 15129
rect 5070 15097 5096 15100
rect 4702 15058 4728 15061
rect 4702 15029 4728 15032
rect 4794 15024 4820 15027
rect 4794 14995 4820 14998
rect 4800 14823 4814 14995
rect 4846 14925 4860 15097
rect 4840 14922 4866 14925
rect 4840 14893 4866 14896
rect 4794 14820 4820 14823
rect 4794 14791 4820 14794
rect 4840 14820 4866 14823
rect 4840 14791 4866 14794
rect 3828 14616 3854 14619
rect 3828 14587 3854 14590
rect 3486 14256 3572 14270
rect 3460 14247 3486 14250
rect 3558 13531 3572 14256
rect 3552 13528 3578 13531
rect 3552 13499 3578 13502
rect 3460 13494 3486 13497
rect 3460 13465 3486 13468
rect 3466 13191 3480 13465
rect 3460 13188 3486 13191
rect 3460 13159 3486 13162
rect 3368 13154 3394 13157
rect 3368 13125 3394 13128
rect 3466 12953 3480 13159
rect 3834 13117 3848 14587
rect 4794 14276 4820 14279
rect 4794 14247 4820 14250
rect 4800 14041 4814 14247
rect 4794 14038 4820 14041
rect 4794 14009 4820 14012
rect 4610 13494 4636 13497
rect 4610 13465 4636 13468
rect 4616 13293 4630 13465
rect 4747 13308 4775 13312
rect 4610 13290 4636 13293
rect 4846 13293 4860 14791
rect 4886 14786 4912 14789
rect 4886 14757 4912 14760
rect 4932 14786 4958 14789
rect 4932 14757 4958 14760
rect 4892 14536 4906 14757
rect 4938 14653 4952 14757
rect 4932 14650 4958 14653
rect 4932 14621 4958 14624
rect 4885 14532 4913 14536
rect 4885 14499 4913 14504
rect 4984 14381 4998 15097
rect 5024 15058 5050 15061
rect 5024 15029 5050 15032
rect 4978 14378 5004 14381
rect 4978 14349 5004 14352
rect 4978 14310 5004 14313
rect 4978 14281 5004 14284
rect 4747 13275 4775 13280
rect 4840 13290 4866 13293
rect 4610 13261 4636 13264
rect 4754 13191 4768 13275
rect 4840 13261 4866 13264
rect 4846 13191 4860 13261
rect 4748 13188 4774 13191
rect 4748 13159 4774 13162
rect 4840 13188 4866 13191
rect 4840 13159 4866 13162
rect 4656 13154 4682 13157
rect 4656 13125 4682 13128
rect 4794 13154 4820 13157
rect 4794 13125 4820 13128
rect 3834 13103 3894 13117
rect 3880 12987 3894 13103
rect 3874 12984 3900 12987
rect 3874 12955 3900 12958
rect 3460 12950 3486 12953
rect 3460 12921 3486 12924
rect 3920 12950 3946 12953
rect 3920 12921 3946 12924
rect 3138 12916 3164 12919
rect 3138 12887 3164 12890
rect 3144 12681 3158 12887
rect 3138 12678 3164 12681
rect 3138 12649 3164 12652
rect 3144 12443 3158 12649
rect 3466 12647 3480 12921
rect 3460 12644 3486 12647
rect 3413 12628 3441 12632
rect 3460 12615 3486 12618
rect 3413 12595 3414 12600
rect 3440 12595 3441 12600
rect 3414 12581 3440 12584
rect 3926 12579 3940 12921
rect 4662 12749 4676 13125
rect 4800 13021 4814 13125
rect 4794 13018 4820 13021
rect 4794 12989 4820 12992
rect 4656 12746 4682 12749
rect 4656 12717 4682 12720
rect 4984 12613 4998 14281
rect 5030 13565 5044 15029
rect 5024 13562 5050 13565
rect 5024 13533 5050 13536
rect 5024 13494 5050 13497
rect 5076 13488 5090 15097
rect 5116 15024 5142 15027
rect 5116 14995 5142 14998
rect 5122 14857 5136 14995
rect 5116 14854 5142 14857
rect 5116 14825 5142 14828
rect 5116 14276 5142 14279
rect 5116 14247 5142 14250
rect 5122 13701 5136 14247
rect 5116 13698 5142 13701
rect 5116 13669 5142 13672
rect 5168 13573 5182 15131
rect 5260 14313 5274 18531
rect 5398 18359 5412 23062
rect 5536 22949 5550 23495
rect 5438 22946 5464 22949
rect 5438 22917 5464 22920
rect 5530 22946 5556 22949
rect 5530 22917 5556 22920
rect 5760 22946 5786 22949
rect 5760 22917 5786 22920
rect 5444 18588 5458 22917
rect 5536 22430 5550 22917
rect 5576 22436 5602 22439
rect 5536 22416 5576 22430
rect 5576 22407 5602 22410
rect 5622 22436 5648 22439
rect 5622 22407 5648 22410
rect 5484 21892 5510 21895
rect 5484 21863 5510 21866
rect 5490 21393 5504 21863
rect 5490 21379 5596 21393
rect 5582 21351 5596 21379
rect 5576 21348 5602 21351
rect 5576 21319 5602 21322
rect 5530 21314 5556 21317
rect 5530 21285 5556 21288
rect 5536 21257 5550 21285
rect 5628 21257 5642 22407
rect 5714 21994 5740 21997
rect 5714 21965 5740 21968
rect 5720 21393 5734 21965
rect 5536 21243 5642 21257
rect 5674 21379 5734 21393
rect 5530 20736 5556 20739
rect 5530 20707 5556 20710
rect 5536 20637 5550 20707
rect 5530 20634 5556 20637
rect 5530 20605 5556 20608
rect 5536 20365 5550 20605
rect 5530 20362 5556 20365
rect 5530 20333 5556 20336
rect 5530 19716 5556 19719
rect 5530 19687 5556 19690
rect 5536 19432 5550 19687
rect 5529 19428 5557 19432
rect 5529 19395 5557 19400
rect 5536 19081 5550 19395
rect 5582 19175 5596 21243
rect 5674 20707 5688 21379
rect 5714 21348 5740 21351
rect 5714 21319 5740 21322
rect 5628 20693 5688 20707
rect 5628 19685 5642 20693
rect 5720 20637 5734 21319
rect 5766 20792 5780 22917
rect 5812 21113 5826 24685
rect 5852 24374 5878 24377
rect 5852 24345 5878 24348
rect 5806 21110 5832 21113
rect 5806 21081 5832 21084
rect 5858 20849 5872 24345
rect 5944 22912 5970 22915
rect 5944 22883 5970 22886
rect 5950 22439 5964 22883
rect 5944 22436 5970 22439
rect 5944 22407 5970 22410
rect 5812 20835 5872 20849
rect 5759 20788 5787 20792
rect 5759 20755 5760 20760
rect 5786 20755 5787 20760
rect 5760 20741 5786 20744
rect 5812 20707 5826 20835
rect 5851 20788 5879 20792
rect 5851 20755 5879 20760
rect 5766 20693 5826 20707
rect 5714 20634 5740 20637
rect 5714 20605 5740 20608
rect 5766 20263 5780 20693
rect 5760 20260 5786 20263
rect 5760 20231 5786 20234
rect 5668 19988 5694 19991
rect 5668 19959 5694 19962
rect 5674 19821 5688 19959
rect 5668 19818 5694 19821
rect 5668 19789 5694 19792
rect 5622 19682 5648 19685
rect 5622 19653 5648 19656
rect 5674 19277 5688 19789
rect 5668 19274 5694 19277
rect 5668 19245 5694 19248
rect 5806 19274 5832 19277
rect 5806 19245 5832 19248
rect 5576 19172 5602 19175
rect 5576 19143 5602 19146
rect 5576 19104 5602 19107
rect 5536 19078 5576 19081
rect 5536 19075 5602 19078
rect 5536 19067 5596 19075
rect 5484 18594 5510 18597
rect 5444 18574 5484 18588
rect 5484 18565 5510 18568
rect 5582 18393 5596 19067
rect 5674 18733 5688 19245
rect 5668 18730 5694 18733
rect 5668 18701 5694 18704
rect 5576 18390 5602 18393
rect 5576 18361 5602 18364
rect 5392 18356 5418 18359
rect 5392 18327 5418 18330
rect 5300 18288 5326 18291
rect 5300 18259 5326 18262
rect 5306 18121 5320 18259
rect 5300 18118 5326 18121
rect 5300 18089 5326 18092
rect 5398 16157 5412 18327
rect 5674 18189 5688 18701
rect 5812 18631 5826 19245
rect 5806 18628 5832 18631
rect 5806 18599 5832 18602
rect 5668 18186 5694 18189
rect 5668 18157 5694 18160
rect 5576 18050 5602 18053
rect 5576 18021 5602 18024
rect 5398 16143 5458 16157
rect 5392 16112 5418 16115
rect 5392 16083 5418 16086
rect 5398 15877 5412 16083
rect 5444 15877 5458 16143
rect 5392 15874 5418 15877
rect 5444 15863 5504 15877
rect 5392 15845 5418 15848
rect 5254 14310 5280 14313
rect 5254 14281 5280 14284
rect 5254 14038 5280 14041
rect 5254 14009 5280 14012
rect 5208 13936 5234 13939
rect 5208 13907 5234 13910
rect 5214 13735 5228 13907
rect 5208 13732 5234 13735
rect 5208 13703 5234 13706
rect 5050 13474 5090 13488
rect 5122 13559 5182 13573
rect 5024 13465 5050 13468
rect 5122 13429 5136 13559
rect 5162 13494 5188 13497
rect 5162 13465 5188 13468
rect 5116 13426 5142 13429
rect 5116 13397 5142 13400
rect 5168 13225 5182 13465
rect 5214 13225 5228 13703
rect 5162 13222 5188 13225
rect 5162 13193 5188 13196
rect 5208 13222 5234 13225
rect 5208 13193 5234 13196
rect 5260 12647 5274 14009
rect 5392 13698 5418 13701
rect 5392 13669 5418 13672
rect 5346 13222 5372 13225
rect 5346 13193 5372 13196
rect 5300 13154 5326 13157
rect 5300 13125 5326 13128
rect 5306 13021 5320 13125
rect 5300 13018 5326 13021
rect 5300 12989 5326 12992
rect 5352 12749 5366 13193
rect 5398 13191 5412 13669
rect 5392 13188 5418 13191
rect 5392 13159 5418 13162
rect 5346 12746 5372 12749
rect 5346 12717 5372 12720
rect 5254 12644 5280 12647
rect 5254 12615 5280 12618
rect 4748 12610 4774 12613
rect 4748 12581 4774 12584
rect 4978 12610 5004 12613
rect 4978 12581 5004 12584
rect 3920 12576 3946 12579
rect 3920 12547 3946 12550
rect 4754 12443 4768 12581
rect 5254 12576 5280 12579
rect 5254 12547 5280 12550
rect 5260 12477 5274 12547
rect 5254 12474 5280 12477
rect 5254 12445 5280 12448
rect 3138 12440 3164 12443
rect 3138 12411 3164 12414
rect 4748 12440 4774 12443
rect 4748 12411 4774 12414
rect 4518 12372 4544 12375
rect 4518 12343 4544 12346
rect 4524 12137 4538 12343
rect 4518 12134 4544 12137
rect 4518 12105 4544 12108
rect 4524 11321 4538 12105
rect 4754 11355 4768 12411
rect 5438 12304 5464 12307
rect 5438 12275 5464 12278
rect 5392 12168 5418 12171
rect 5392 12139 5418 12142
rect 4840 12066 4866 12069
rect 4840 12037 4866 12040
rect 4846 11933 4860 12037
rect 5398 12020 5412 12139
rect 5391 12016 5419 12020
rect 5391 11983 5419 11988
rect 5398 11933 5412 11983
rect 5444 11933 5458 12275
rect 4840 11930 4866 11933
rect 4840 11901 4866 11904
rect 5392 11930 5418 11933
rect 5392 11901 5418 11904
rect 5438 11930 5464 11933
rect 5438 11901 5464 11904
rect 5490 11831 5504 15863
rect 5582 13117 5596 18021
rect 5674 17543 5688 18157
rect 5760 17880 5786 17883
rect 5760 17851 5786 17854
rect 5766 17543 5780 17851
rect 5668 17540 5694 17543
rect 5668 17511 5694 17514
rect 5760 17540 5786 17543
rect 5760 17511 5786 17514
rect 5674 17101 5688 17511
rect 5766 17305 5780 17511
rect 5858 17509 5872 20755
rect 5996 18053 6010 28731
rect 6680 28731 6706 28734
rect 6587 28711 6588 28716
rect 6614 28711 6615 28716
rect 6588 28697 6614 28700
rect 6686 28423 6700 28731
rect 6680 28420 6706 28423
rect 6680 28391 6706 28394
rect 6686 27641 6700 28391
rect 6680 27638 6706 27641
rect 6680 27609 6706 27612
rect 6358 27536 6384 27539
rect 6358 27507 6384 27510
rect 6266 27366 6292 27369
rect 6266 27337 6292 27340
rect 6036 27332 6062 27335
rect 6036 27303 6062 27306
rect 6042 27165 6056 27303
rect 6272 27165 6286 27337
rect 6036 27162 6062 27165
rect 6036 27133 6062 27136
rect 6266 27162 6292 27165
rect 6266 27133 6292 27136
rect 6220 27094 6246 27097
rect 6220 27065 6246 27068
rect 6226 26621 6240 27065
rect 6364 27063 6378 27507
rect 6732 27437 6746 29207
rect 6962 29069 6976 29241
rect 6956 29066 6982 29069
rect 6956 29037 6982 29040
rect 6818 28964 6844 28967
rect 6818 28935 6844 28938
rect 6864 28964 6890 28967
rect 6864 28935 6890 28938
rect 6824 28797 6838 28935
rect 6818 28794 6844 28797
rect 6818 28765 6844 28768
rect 6818 28726 6844 28729
rect 6818 28697 6844 28700
rect 6772 28420 6798 28423
rect 6772 28391 6798 28394
rect 6824 28397 6838 28697
rect 6870 28491 6884 28935
rect 6956 28794 6982 28797
rect 6956 28765 6982 28768
rect 6962 28729 6976 28765
rect 6956 28726 6982 28729
rect 6956 28697 6982 28700
rect 6864 28488 6890 28491
rect 6864 28459 6890 28462
rect 6778 27709 6792 28391
rect 6824 28383 6884 28397
rect 6772 27706 6798 27709
rect 6772 27677 6798 27680
rect 6726 27434 6752 27437
rect 6726 27405 6752 27408
rect 6732 27097 6746 27405
rect 6772 27264 6798 27267
rect 6772 27235 6798 27238
rect 6778 27131 6792 27235
rect 6772 27128 6798 27131
rect 6772 27099 6798 27102
rect 6726 27094 6752 27097
rect 6726 27065 6752 27068
rect 6358 27060 6384 27063
rect 6358 27031 6384 27034
rect 6634 26788 6660 26791
rect 6634 26759 6660 26762
rect 6640 26621 6654 26759
rect 6220 26618 6246 26621
rect 6220 26589 6246 26592
rect 6634 26618 6660 26621
rect 6634 26589 6660 26592
rect 6220 26550 6246 26553
rect 6220 26521 6246 26524
rect 6226 26349 6240 26521
rect 6220 26346 6246 26349
rect 6220 26317 6246 26320
rect 6778 26213 6792 27099
rect 6870 26791 6884 28383
rect 6962 27675 6976 28697
rect 6956 27672 6982 27675
rect 6956 27643 6982 27646
rect 6956 27604 6982 27607
rect 6956 27575 6982 27578
rect 6962 27403 6976 27575
rect 6956 27400 6982 27403
rect 6956 27371 6982 27374
rect 6910 26856 6936 26859
rect 6910 26827 6936 26830
rect 6962 26833 6976 27371
rect 7054 27267 7068 29275
rect 8710 29273 8724 29445
rect 10274 29307 10288 29547
rect 10360 29508 10386 29511
rect 10360 29479 10386 29482
rect 10498 29508 10524 29511
rect 10498 29479 10524 29482
rect 11372 29508 11398 29511
rect 11372 29479 11398 29482
rect 12292 29508 12318 29511
rect 12292 29479 12318 29482
rect 10268 29304 10294 29307
rect 10268 29275 10294 29278
rect 8704 29270 8730 29273
rect 8704 29241 8730 29244
rect 8796 29270 8822 29273
rect 8796 29241 8822 29244
rect 9026 29270 9052 29273
rect 9026 29241 9052 29244
rect 10314 29270 10340 29273
rect 10314 29241 10340 29244
rect 8060 29168 8086 29171
rect 8060 29139 8086 29142
rect 8066 28967 8080 29139
rect 8658 29032 8684 29035
rect 8658 29003 8684 29006
rect 7462 28964 7488 28967
rect 7330 28938 7462 28941
rect 7330 28935 7488 28938
rect 7508 28964 7534 28967
rect 7508 28935 7534 28938
rect 8060 28964 8086 28967
rect 8060 28935 8086 28938
rect 8428 28964 8454 28967
rect 8428 28935 8454 28938
rect 7330 28933 7482 28935
rect 7324 28930 7482 28933
rect 7350 28927 7482 28930
rect 7324 28901 7350 28904
rect 7376 27675 7390 28927
rect 7514 28763 7528 28935
rect 7508 28760 7534 28763
rect 7508 28731 7534 28734
rect 7692 28726 7718 28729
rect 7692 28697 7718 28700
rect 7370 27672 7396 27675
rect 7370 27643 7396 27646
rect 7186 27638 7212 27641
rect 7186 27609 7212 27612
rect 7048 27264 7074 27267
rect 7048 27235 7074 27238
rect 6864 26788 6890 26791
rect 6864 26759 6890 26762
rect 6870 26519 6884 26759
rect 6864 26516 6890 26519
rect 6864 26487 6890 26490
rect 6772 26210 6798 26213
rect 6772 26181 6798 26184
rect 6082 25904 6108 25907
rect 6082 25875 6108 25878
rect 6634 25904 6660 25907
rect 6634 25875 6660 25878
rect 6088 24921 6102 25875
rect 6174 25632 6200 25635
rect 6174 25603 6200 25606
rect 6180 24921 6194 25603
rect 6640 25465 6654 25875
rect 6778 25499 6792 26181
rect 6916 26077 6930 26827
rect 6962 26825 7022 26833
rect 6962 26822 7028 26825
rect 6962 26819 7002 26822
rect 6962 26553 6976 26819
rect 7002 26793 7028 26796
rect 7002 26754 7028 26757
rect 7002 26725 7028 26728
rect 6956 26550 6982 26553
rect 6956 26521 6982 26524
rect 6910 26074 6936 26077
rect 6910 26045 6936 26048
rect 7008 25975 7022 26725
rect 7192 26621 7206 27609
rect 7376 27369 7390 27643
rect 7698 27607 7712 28697
rect 7600 27604 7626 27607
rect 7600 27575 7626 27578
rect 7692 27604 7718 27607
rect 7692 27575 7718 27578
rect 7370 27366 7396 27369
rect 7370 27337 7396 27340
rect 7606 27335 7620 27575
rect 7646 27536 7672 27539
rect 7646 27507 7672 27510
rect 7652 27369 7666 27507
rect 7646 27366 7672 27369
rect 7646 27337 7672 27340
rect 7508 27332 7534 27335
rect 7508 27303 7534 27306
rect 7600 27332 7626 27335
rect 7600 27303 7626 27306
rect 7416 27264 7442 27267
rect 7416 27235 7442 27238
rect 7422 27097 7436 27235
rect 7416 27094 7442 27097
rect 7416 27065 7442 27068
rect 7416 26992 7442 26995
rect 7416 26963 7442 26966
rect 7278 26720 7304 26723
rect 7278 26691 7304 26694
rect 7186 26618 7212 26621
rect 7186 26589 7212 26592
rect 7192 26553 7206 26589
rect 7284 26553 7298 26691
rect 7186 26550 7212 26553
rect 7186 26521 7212 26524
rect 7278 26550 7304 26553
rect 7278 26521 7304 26524
rect 7232 26176 7258 26179
rect 7232 26147 7258 26150
rect 7048 26006 7074 26009
rect 7048 25977 7074 25980
rect 7002 25972 7028 25975
rect 7002 25943 7028 25946
rect 7054 25805 7068 25977
rect 7048 25802 7074 25805
rect 7048 25773 7074 25776
rect 6772 25496 6798 25499
rect 6772 25467 6798 25470
rect 6634 25462 6660 25465
rect 6634 25433 6660 25436
rect 6358 25088 6384 25091
rect 6358 25059 6384 25062
rect 6082 24918 6108 24921
rect 6082 24889 6108 24892
rect 6174 24918 6200 24921
rect 6174 24889 6200 24892
rect 6220 24612 6246 24615
rect 6220 24583 6246 24586
rect 6036 23728 6062 23731
rect 6036 23699 6062 23702
rect 6042 23561 6056 23699
rect 6036 23558 6062 23561
rect 6036 23529 6062 23532
rect 6226 22481 6240 24583
rect 6364 23867 6378 25059
rect 6542 24884 6568 24887
rect 6542 24855 6568 24858
rect 6496 24850 6522 24853
rect 6496 24821 6522 24824
rect 6404 24816 6430 24819
rect 6404 24787 6430 24790
rect 6358 23864 6384 23867
rect 6358 23835 6384 23838
rect 6358 23728 6384 23731
rect 6358 23699 6384 23702
rect 6364 23527 6378 23699
rect 6410 23595 6424 24787
rect 6502 24275 6516 24821
rect 6548 24717 6562 24855
rect 6542 24714 6568 24717
rect 6542 24685 6568 24688
rect 6956 24646 6982 24649
rect 6956 24617 6982 24620
rect 6910 24340 6936 24343
rect 6910 24311 6936 24314
rect 6496 24272 6522 24275
rect 6496 24243 6522 24246
rect 6450 23830 6476 23833
rect 6450 23801 6476 23804
rect 6404 23592 6430 23595
rect 6404 23563 6430 23566
rect 6358 23524 6384 23527
rect 6358 23495 6384 23498
rect 6266 23456 6292 23459
rect 6266 23427 6292 23430
rect 6312 23456 6338 23459
rect 6312 23427 6338 23430
rect 6272 23323 6286 23427
rect 6266 23320 6292 23323
rect 6266 23291 6292 23294
rect 6318 23255 6332 23427
rect 6404 23286 6430 23289
rect 6404 23257 6430 23260
rect 6312 23252 6338 23255
rect 6312 23223 6338 23226
rect 6410 22541 6424 23257
rect 6456 23085 6470 23801
rect 6450 23082 6476 23085
rect 6450 23053 6476 23056
rect 6404 22538 6430 22541
rect 6404 22509 6430 22512
rect 6226 22467 6424 22481
rect 6358 20736 6384 20739
rect 6358 20707 6384 20710
rect 6364 20603 6378 20707
rect 6358 20600 6384 20603
rect 6358 20571 6384 20574
rect 6174 20532 6200 20535
rect 6174 20503 6200 20506
rect 6082 20260 6108 20263
rect 6082 20231 6108 20234
rect 6036 18458 6062 18461
rect 6036 18429 6062 18432
rect 6042 18189 6056 18429
rect 6036 18186 6062 18189
rect 6036 18157 6062 18160
rect 5990 18050 6016 18053
rect 5990 18021 6016 18024
rect 5852 17506 5878 17509
rect 5852 17477 5878 17480
rect 5760 17302 5786 17305
rect 5760 17273 5786 17276
rect 5668 17098 5694 17101
rect 5668 17069 5694 17072
rect 5674 16455 5688 17069
rect 5766 16999 5780 17273
rect 5760 16996 5786 16999
rect 5760 16967 5786 16970
rect 5668 16452 5694 16455
rect 5694 16432 5734 16446
rect 5668 16423 5694 16426
rect 5622 16418 5648 16421
rect 5622 16389 5648 16392
rect 5628 15741 5642 16389
rect 5720 15911 5734 16432
rect 5714 15908 5740 15911
rect 5714 15879 5740 15882
rect 5760 15908 5786 15911
rect 5760 15879 5786 15882
rect 5622 15738 5648 15741
rect 5622 15709 5648 15712
rect 5628 15367 5642 15709
rect 5668 15670 5694 15673
rect 5668 15641 5694 15644
rect 5622 15364 5648 15367
rect 5622 15335 5648 15338
rect 5674 13117 5688 15641
rect 5720 15469 5734 15879
rect 5766 15673 5780 15879
rect 5760 15670 5786 15673
rect 5760 15641 5786 15644
rect 5714 15466 5740 15469
rect 5714 15437 5740 15440
rect 5720 14313 5734 15437
rect 5858 15333 5872 17477
rect 6088 16999 6102 20231
rect 6180 19991 6194 20503
rect 6410 20195 6424 22467
rect 6502 22424 6516 24243
rect 6916 24105 6930 24311
rect 6910 24102 6936 24105
rect 6910 24073 6936 24076
rect 6916 23833 6930 24073
rect 6962 24037 6976 24617
rect 7054 24377 7068 25773
rect 7238 25737 7252 26147
rect 7232 25734 7258 25737
rect 7232 25705 7258 25708
rect 7048 24374 7074 24377
rect 7048 24345 7074 24348
rect 7054 24139 7068 24345
rect 7048 24136 7074 24139
rect 7048 24107 7074 24110
rect 6956 24034 6982 24037
rect 6956 24005 6982 24008
rect 6955 23984 6983 23988
rect 6955 23951 6983 23956
rect 6962 23867 6976 23951
rect 6956 23864 6982 23867
rect 6956 23835 6982 23838
rect 6818 23830 6844 23833
rect 6818 23801 6844 23804
rect 6910 23830 6936 23833
rect 6910 23801 6936 23804
rect 6588 23796 6614 23799
rect 6588 23767 6614 23770
rect 6495 22420 6523 22424
rect 6495 22387 6523 22392
rect 6450 21892 6476 21895
rect 6450 21863 6476 21866
rect 6456 21725 6470 21863
rect 6542 21824 6568 21827
rect 6542 21795 6568 21798
rect 6450 21722 6476 21725
rect 6450 21693 6476 21696
rect 6548 21657 6562 21795
rect 6496 21654 6522 21657
rect 6496 21625 6522 21628
rect 6542 21654 6568 21657
rect 6542 21625 6568 21628
rect 6502 21181 6516 21625
rect 6496 21178 6522 21181
rect 6496 21149 6522 21152
rect 6594 21147 6608 23767
rect 6634 23320 6660 23323
rect 6634 23291 6660 23294
rect 6640 23051 6654 23291
rect 6726 23286 6752 23289
rect 6726 23257 6752 23260
rect 6732 23187 6746 23257
rect 6726 23184 6752 23187
rect 6726 23155 6752 23158
rect 6634 23048 6660 23051
rect 6634 23019 6660 23022
rect 6640 21929 6654 23019
rect 6634 21926 6660 21929
rect 6660 21906 6700 21920
rect 6634 21897 6660 21900
rect 6634 21858 6660 21861
rect 6634 21829 6660 21832
rect 6640 21453 6654 21829
rect 6634 21450 6660 21453
rect 6634 21421 6660 21424
rect 6686 21172 6700 21906
rect 6732 21895 6746 23155
rect 6726 21892 6752 21895
rect 6726 21863 6752 21866
rect 6640 21158 6700 21172
rect 6588 21144 6614 21147
rect 6588 21115 6614 21118
rect 6542 21110 6568 21113
rect 6542 21081 6568 21084
rect 6496 20566 6522 20569
rect 6496 20537 6522 20540
rect 6404 20192 6430 20195
rect 6404 20163 6430 20166
rect 6410 20059 6424 20163
rect 6404 20056 6430 20059
rect 6404 20027 6430 20030
rect 6502 20025 6516 20537
rect 6548 20365 6562 21081
rect 6640 21053 6654 21158
rect 6680 21110 6706 21113
rect 6680 21081 6706 21084
rect 6594 21039 6654 21053
rect 6542 20362 6568 20365
rect 6542 20333 6568 20336
rect 6496 20022 6522 20025
rect 6496 19993 6522 19996
rect 6174 19988 6200 19991
rect 6174 19959 6200 19962
rect 6594 19812 6608 21039
rect 6686 20909 6700 21081
rect 6680 20906 6706 20909
rect 6680 20877 6706 20880
rect 6732 20849 6746 21863
rect 6772 21144 6798 21147
rect 6824 21132 6838 23801
rect 6772 21115 6798 21118
rect 6817 21128 6845 21132
rect 6502 19798 6608 19812
rect 6640 20835 6746 20849
rect 6404 19648 6430 19651
rect 6404 19619 6430 19622
rect 6410 18937 6424 19619
rect 6502 18971 6516 19798
rect 6542 19104 6568 19107
rect 6542 19075 6568 19078
rect 6548 18971 6562 19075
rect 6496 18968 6522 18971
rect 6496 18939 6522 18942
rect 6542 18968 6568 18971
rect 6542 18939 6568 18942
rect 6640 18937 6654 20835
rect 6726 20804 6752 20807
rect 6726 20775 6752 20778
rect 6404 18934 6430 18937
rect 6404 18905 6430 18908
rect 6634 18934 6660 18937
rect 6634 18905 6660 18908
rect 6266 18560 6292 18563
rect 6266 18531 6292 18534
rect 6272 18461 6286 18531
rect 6266 18458 6292 18461
rect 6266 18429 6292 18432
rect 6174 18390 6200 18393
rect 6174 18361 6200 18364
rect 6180 17883 6194 18361
rect 6732 18087 6746 20775
rect 6778 18155 6792 21115
rect 6817 21095 6818 21100
rect 6844 21095 6845 21100
rect 6818 21081 6844 21084
rect 6824 20807 6838 21081
rect 6962 20841 6976 23835
rect 7054 23833 7068 24107
rect 7048 23830 7074 23833
rect 7048 23801 7074 23804
rect 7002 22232 7028 22235
rect 7002 22203 7028 22206
rect 6956 20838 6982 20841
rect 6956 20809 6982 20812
rect 6818 20804 6844 20807
rect 6818 20775 6844 20778
rect 7008 20569 7022 22203
rect 7238 21691 7252 25705
rect 7422 25431 7436 26963
rect 7514 26859 7528 27303
rect 7600 27060 7626 27063
rect 7560 27034 7600 27037
rect 7560 27031 7626 27034
rect 7560 27023 7620 27031
rect 7508 26856 7534 26859
rect 7508 26827 7534 26830
rect 7514 26349 7528 26827
rect 7560 26791 7574 27023
rect 7698 26825 7712 27575
rect 7738 27570 7764 27573
rect 7738 27541 7764 27544
rect 7744 27165 7758 27541
rect 7738 27162 7764 27165
rect 7738 27133 7764 27136
rect 7692 26822 7718 26825
rect 7692 26793 7718 26796
rect 7554 26788 7580 26791
rect 7554 26759 7580 26762
rect 7560 26621 7574 26759
rect 7554 26618 7580 26621
rect 7554 26589 7580 26592
rect 7698 26587 7712 26793
rect 7692 26584 7718 26587
rect 7692 26555 7718 26558
rect 7508 26346 7534 26349
rect 7508 26317 7534 26320
rect 7508 26210 7534 26213
rect 7508 26181 7534 26184
rect 7514 26043 7528 26181
rect 7554 26176 7580 26179
rect 7554 26147 7580 26150
rect 7508 26040 7534 26043
rect 7508 26011 7534 26014
rect 7560 26009 7574 26147
rect 7554 26006 7580 26009
rect 7554 25977 7580 25980
rect 7554 25802 7580 25805
rect 7554 25773 7580 25776
rect 7560 25533 7574 25773
rect 7744 25703 7758 27133
rect 7738 25700 7764 25703
rect 7738 25671 7764 25674
rect 7744 25537 7758 25671
rect 7554 25530 7580 25533
rect 7744 25523 7850 25537
rect 7554 25501 7580 25504
rect 7416 25428 7442 25431
rect 7416 25399 7442 25402
rect 7324 23830 7350 23833
rect 7324 23801 7350 23804
rect 7330 22745 7344 23801
rect 7324 22742 7350 22745
rect 7350 22722 7390 22736
rect 7324 22713 7350 22716
rect 7278 22708 7304 22711
rect 7278 22679 7304 22682
rect 7284 22439 7298 22679
rect 7376 22473 7390 22722
rect 7370 22470 7396 22473
rect 7370 22441 7396 22444
rect 7278 22436 7304 22439
rect 7278 22407 7304 22410
rect 7376 22201 7390 22441
rect 7370 22198 7396 22201
rect 7370 22169 7396 22172
rect 7232 21688 7258 21691
rect 7232 21659 7258 21662
rect 7238 21147 7252 21659
rect 7278 21620 7304 21623
rect 7278 21591 7304 21594
rect 7284 21283 7298 21591
rect 7278 21280 7304 21283
rect 7278 21251 7304 21254
rect 7232 21144 7258 21147
rect 7232 21115 7258 21118
rect 7238 20739 7252 21115
rect 7284 21079 7298 21251
rect 7278 21076 7304 21079
rect 7278 21047 7304 21050
rect 7232 20736 7258 20739
rect 7232 20707 7258 20710
rect 7002 20566 7028 20569
rect 7002 20537 7028 20540
rect 7008 19704 7022 20537
rect 7048 20192 7074 20195
rect 7048 20163 7074 20166
rect 7001 19700 7029 19704
rect 7001 19667 7029 19672
rect 6818 19138 6844 19141
rect 6818 19109 6844 19112
rect 6910 19138 6936 19141
rect 6910 19109 6936 19112
rect 6824 19005 6838 19109
rect 6818 19002 6844 19005
rect 6818 18973 6844 18976
rect 6916 18189 6930 19109
rect 6956 18900 6982 18903
rect 6956 18871 6982 18874
rect 6962 18393 6976 18871
rect 7008 18393 7022 19667
rect 6956 18390 6982 18393
rect 6956 18361 6982 18364
rect 7002 18390 7028 18393
rect 7002 18361 7028 18364
rect 6956 18288 6982 18291
rect 6956 18259 6982 18262
rect 6910 18186 6936 18189
rect 6910 18157 6936 18160
rect 6772 18152 6798 18155
rect 6772 18123 6798 18126
rect 6680 18084 6706 18087
rect 6680 18055 6706 18058
rect 6726 18084 6752 18087
rect 6726 18055 6752 18058
rect 6174 17880 6200 17883
rect 6174 17851 6200 17854
rect 6686 17101 6700 18055
rect 6778 18053 6792 18123
rect 6864 18084 6890 18087
rect 6864 18055 6890 18058
rect 6772 18050 6798 18053
rect 6772 18021 6798 18024
rect 6818 18050 6844 18053
rect 6818 18021 6844 18024
rect 6824 17645 6838 18021
rect 6818 17642 6844 17645
rect 6818 17613 6844 17616
rect 6680 17098 6706 17101
rect 6680 17069 6706 17072
rect 6082 16996 6108 16999
rect 6082 16967 6108 16970
rect 6312 16656 6338 16659
rect 6312 16627 6338 16630
rect 6318 16455 6332 16627
rect 6772 16554 6798 16557
rect 6772 16525 6798 16528
rect 6312 16452 6338 16455
rect 6778 16440 6792 16525
rect 6312 16423 6338 16426
rect 6771 16436 6799 16440
rect 5990 16418 6016 16421
rect 5990 16389 6016 16392
rect 5996 16304 6010 16389
rect 5989 16300 6017 16304
rect 5989 16267 6017 16272
rect 6318 16217 6332 16423
rect 6771 16403 6799 16408
rect 6726 16384 6752 16387
rect 6726 16355 6752 16358
rect 6732 16285 6746 16355
rect 6726 16282 6752 16285
rect 6726 16253 6752 16256
rect 6778 16217 6792 16403
rect 6266 16214 6292 16217
rect 6266 16185 6292 16188
rect 6312 16214 6338 16217
rect 6312 16185 6338 16188
rect 6772 16214 6798 16217
rect 6772 16185 6798 16188
rect 6272 16013 6286 16185
rect 6634 16112 6660 16115
rect 6634 16083 6660 16086
rect 6266 16010 6292 16013
rect 6266 15981 6292 15984
rect 5990 15364 6016 15367
rect 5990 15335 6016 15338
rect 5852 15330 5878 15333
rect 5852 15301 5878 15304
rect 5944 15194 5970 15197
rect 5944 15165 5970 15168
rect 5898 14820 5924 14823
rect 5898 14791 5924 14794
rect 5904 14585 5918 14791
rect 5950 14755 5964 15165
rect 5996 14814 6010 15335
rect 6640 15129 6654 16083
rect 6772 15296 6798 15299
rect 6772 15267 6798 15270
rect 6778 15129 6792 15267
rect 6870 15163 6884 18055
rect 6962 17849 6976 18259
rect 7054 17857 7068 20163
rect 7284 19481 7298 21047
rect 7422 19481 7436 25399
rect 7784 24918 7810 24921
rect 7784 24889 7810 24892
rect 7738 24578 7764 24581
rect 7738 24549 7764 24552
rect 7744 24445 7758 24549
rect 7738 24442 7764 24445
rect 7738 24413 7764 24416
rect 7554 24374 7580 24377
rect 7554 24345 7580 24348
rect 7560 24037 7574 24345
rect 7554 24034 7580 24037
rect 7554 24005 7580 24008
rect 7560 22821 7574 24005
rect 7514 22807 7574 22821
rect 7462 22402 7488 22405
rect 7462 22373 7488 22376
rect 7468 22099 7482 22373
rect 7462 22096 7488 22099
rect 7462 22067 7488 22070
rect 7468 21283 7482 22067
rect 7462 21280 7488 21283
rect 7462 21251 7488 21254
rect 7468 20841 7482 21251
rect 7514 21147 7528 22807
rect 7554 22742 7580 22745
rect 7554 22713 7580 22716
rect 7508 21144 7534 21147
rect 7508 21115 7534 21118
rect 7514 20909 7528 21115
rect 7508 20906 7534 20909
rect 7508 20877 7534 20880
rect 7462 20838 7488 20841
rect 7462 20809 7488 20812
rect 7278 19478 7304 19481
rect 7278 19449 7304 19452
rect 7416 19478 7442 19481
rect 7416 19449 7442 19452
rect 7284 19209 7298 19449
rect 7278 19206 7304 19209
rect 7278 19177 7304 19180
rect 7284 18937 7298 19177
rect 7422 19141 7436 19449
rect 7416 19138 7442 19141
rect 7416 19109 7442 19112
rect 7422 18937 7436 19109
rect 7514 18971 7528 20877
rect 7560 20807 7574 22713
rect 7646 22402 7672 22405
rect 7646 22373 7672 22376
rect 7652 22345 7666 22373
rect 7606 22331 7666 22345
rect 7606 21657 7620 22331
rect 7600 21654 7626 21657
rect 7600 21625 7626 21628
rect 7554 20804 7580 20807
rect 7554 20775 7580 20778
rect 7560 19515 7574 20775
rect 7606 20603 7620 21625
rect 7646 21552 7672 21555
rect 7646 21523 7672 21526
rect 7652 21453 7666 21523
rect 7646 21450 7672 21453
rect 7646 21421 7672 21424
rect 7790 20707 7804 24889
rect 7836 23705 7850 25523
rect 8066 25397 8080 28935
rect 8152 28930 8178 28933
rect 8152 28901 8178 28904
rect 8158 28729 8172 28901
rect 8434 28797 8448 28935
rect 8382 28794 8408 28797
rect 8382 28765 8408 28768
rect 8428 28794 8454 28797
rect 8428 28765 8454 28768
rect 8388 28729 8402 28765
rect 8664 28763 8678 29003
rect 8658 28760 8684 28763
rect 8658 28731 8684 28734
rect 8152 28726 8178 28729
rect 8152 28697 8178 28700
rect 8382 28726 8408 28729
rect 8382 28697 8408 28700
rect 8290 28624 8316 28627
rect 8290 28595 8316 28598
rect 8296 28389 8310 28595
rect 8290 28386 8316 28389
rect 8290 28357 8316 28360
rect 8664 28083 8678 28731
rect 8710 28389 8724 29241
rect 8802 29009 8816 29241
rect 8934 29168 8960 29171
rect 8934 29139 8960 29142
rect 8888 29032 8914 29035
rect 8802 29006 8888 29009
rect 8802 29003 8914 29006
rect 8802 28995 8908 29003
rect 8802 28729 8816 28995
rect 8940 28967 8954 29139
rect 8934 28964 8960 28967
rect 8934 28935 8960 28938
rect 8796 28726 8822 28729
rect 8796 28697 8822 28700
rect 8704 28386 8730 28389
rect 8704 28357 8730 28360
rect 8940 28185 8954 28935
rect 9032 28729 9046 29241
rect 10320 29213 10334 29241
rect 10228 29199 10334 29213
rect 9302 28930 9328 28933
rect 9302 28901 9328 28904
rect 9026 28726 9052 28729
rect 9026 28697 9052 28700
rect 8980 28692 9006 28695
rect 8980 28663 9006 28666
rect 8986 28253 9000 28663
rect 9118 28352 9144 28355
rect 9118 28323 9144 28326
rect 8980 28250 9006 28253
rect 8980 28221 9006 28224
rect 9124 28185 9138 28323
rect 9308 28219 9322 28901
rect 9348 28692 9374 28695
rect 9348 28663 9374 28666
rect 9302 28216 9328 28219
rect 9302 28187 9328 28190
rect 8750 28182 8776 28185
rect 8750 28153 8776 28156
rect 8934 28182 8960 28185
rect 8934 28153 8960 28156
rect 9118 28182 9144 28185
rect 9118 28153 9144 28156
rect 8658 28080 8684 28083
rect 8658 28051 8684 28054
rect 8664 27675 8678 28051
rect 8658 27672 8684 27675
rect 8658 27643 8684 27646
rect 8664 27335 8678 27643
rect 8756 27403 8770 28153
rect 8750 27400 8776 27403
rect 8750 27371 8776 27374
rect 8658 27332 8684 27335
rect 8618 27312 8658 27326
rect 8152 27264 8178 27267
rect 8152 27235 8178 27238
rect 8158 27131 8172 27235
rect 8152 27128 8178 27131
rect 8152 27099 8178 27102
rect 8198 27128 8224 27131
rect 8198 27099 8224 27102
rect 8204 26825 8218 27099
rect 8336 26992 8362 26995
rect 8336 26963 8362 26966
rect 8198 26822 8224 26825
rect 8198 26793 8224 26796
rect 8342 26281 8356 26963
rect 8618 26791 8632 27312
rect 8658 27303 8684 27306
rect 8750 27298 8776 27301
rect 8750 27269 8776 27272
rect 8756 27097 8770 27269
rect 8750 27094 8776 27097
rect 8750 27065 8776 27068
rect 8658 26992 8684 26995
rect 8658 26963 8684 26966
rect 8664 26825 8678 26963
rect 8658 26822 8684 26825
rect 8658 26793 8684 26796
rect 8612 26788 8638 26791
rect 8612 26759 8638 26762
rect 8934 26754 8960 26757
rect 8934 26725 8960 26728
rect 8474 26720 8500 26723
rect 8474 26691 8500 26694
rect 8566 26720 8592 26723
rect 8566 26691 8592 26694
rect 8336 26278 8362 26281
rect 8336 26249 8362 26252
rect 8480 26247 8494 26691
rect 8572 26349 8586 26691
rect 8566 26346 8592 26349
rect 8566 26317 8592 26320
rect 8428 26244 8454 26247
rect 8428 26215 8454 26218
rect 8474 26244 8500 26247
rect 8474 26215 8500 26218
rect 8244 26210 8270 26213
rect 8244 26181 8270 26184
rect 8250 25907 8264 26181
rect 8434 25975 8448 26215
rect 8704 26210 8730 26213
rect 8704 26181 8730 26184
rect 8710 26009 8724 26181
rect 8940 26179 8954 26725
rect 9072 26448 9098 26451
rect 9072 26419 9098 26422
rect 8934 26176 8960 26179
rect 8934 26147 8960 26150
rect 8704 26006 8730 26009
rect 8704 25977 8730 25980
rect 8428 25972 8454 25975
rect 8428 25943 8454 25946
rect 8842 25972 8868 25975
rect 8842 25943 8868 25946
rect 8244 25904 8270 25907
rect 8244 25875 8270 25878
rect 8250 25635 8264 25875
rect 8520 25700 8546 25703
rect 8520 25671 8546 25674
rect 8106 25632 8132 25635
rect 8106 25603 8132 25606
rect 8244 25632 8270 25635
rect 8244 25603 8270 25606
rect 8060 25394 8086 25397
rect 8060 25365 8086 25368
rect 7922 24612 7948 24615
rect 7922 24583 7948 24586
rect 7876 24578 7902 24581
rect 7876 24549 7902 24552
rect 7882 23799 7896 24549
rect 7928 24453 7942 24583
rect 8060 24544 8086 24547
rect 8060 24515 8086 24518
rect 7928 24445 8034 24453
rect 7928 24442 8040 24445
rect 7928 24439 8014 24442
rect 7876 23796 7902 23799
rect 7876 23767 7902 23770
rect 7836 23691 7896 23705
rect 7790 20693 7850 20707
rect 7600 20600 7626 20603
rect 7600 20571 7626 20574
rect 7836 20569 7850 20693
rect 7692 20566 7718 20569
rect 7692 20537 7718 20540
rect 7784 20566 7810 20569
rect 7784 20537 7810 20540
rect 7830 20566 7856 20569
rect 7830 20537 7856 20540
rect 7698 20501 7712 20537
rect 7646 20498 7672 20501
rect 7646 20469 7672 20472
rect 7692 20498 7718 20501
rect 7692 20469 7718 20472
rect 7554 19512 7580 19515
rect 7554 19483 7580 19486
rect 7508 18968 7534 18971
rect 7508 18939 7534 18942
rect 7278 18934 7304 18937
rect 7278 18905 7304 18908
rect 7416 18934 7442 18937
rect 7416 18905 7442 18908
rect 7094 18390 7120 18393
rect 7094 18361 7120 18364
rect 7008 17849 7068 17857
rect 6956 17846 6982 17849
rect 6956 17817 6982 17820
rect 7002 17846 7068 17849
rect 7028 17843 7068 17846
rect 7002 17817 7028 17820
rect 6962 17305 6976 17817
rect 6956 17302 6982 17305
rect 6956 17273 6982 17276
rect 7008 15877 7022 17817
rect 7048 16996 7074 16999
rect 7048 16967 7074 16970
rect 6962 15863 7022 15877
rect 6864 15160 6890 15163
rect 6864 15131 6890 15134
rect 6450 15126 6476 15129
rect 6450 15097 6476 15100
rect 6634 15126 6660 15129
rect 6634 15097 6660 15100
rect 6772 15126 6798 15129
rect 6772 15097 6798 15100
rect 6910 15126 6936 15129
rect 6910 15097 6936 15100
rect 6404 15024 6430 15027
rect 6404 14995 6430 14998
rect 6036 14820 6062 14823
rect 5996 14800 6036 14814
rect 6036 14791 6062 14794
rect 5944 14752 5970 14755
rect 5944 14723 5970 14726
rect 6042 14604 6056 14791
rect 6128 14786 6154 14789
rect 6128 14757 6154 14760
rect 6035 14600 6063 14604
rect 5898 14582 5924 14585
rect 6035 14567 6063 14572
rect 5898 14553 5924 14556
rect 5714 14310 5740 14313
rect 5714 14281 5740 14284
rect 5720 13735 5734 14281
rect 6042 14279 6056 14567
rect 6036 14276 6062 14279
rect 6036 14247 6062 14250
rect 5714 13732 5740 13735
rect 5714 13703 5740 13706
rect 5536 13103 5596 13117
rect 5628 13103 5688 13117
rect 5536 12069 5550 13103
rect 5628 13021 5642 13103
rect 5622 13018 5648 13021
rect 5622 12989 5648 12992
rect 5628 12477 5642 12989
rect 5622 12474 5648 12477
rect 5622 12445 5648 12448
rect 5944 12474 5970 12477
rect 5944 12445 5970 12448
rect 5950 12103 5964 12445
rect 5852 12100 5878 12103
rect 5944 12100 5970 12103
rect 5878 12074 5918 12077
rect 5852 12071 5918 12074
rect 5944 12071 5970 12074
rect 5530 12066 5556 12069
rect 5530 12037 5556 12040
rect 5668 12066 5694 12069
rect 5858 12063 5918 12071
rect 5668 12037 5694 12040
rect 5346 11828 5372 11831
rect 5346 11799 5372 11802
rect 5484 11828 5510 11831
rect 5484 11799 5510 11802
rect 4748 11352 4774 11355
rect 4748 11323 4774 11326
rect 4518 11318 4544 11321
rect 4518 11289 4544 11292
rect 4754 10811 4768 11323
rect 5352 11049 5366 11799
rect 5622 11284 5648 11287
rect 5622 11255 5648 11258
rect 5530 11216 5556 11219
rect 5530 11187 5556 11190
rect 5346 11046 5372 11049
rect 5346 11017 5372 11020
rect 5116 10944 5142 10947
rect 5116 10915 5142 10918
rect 5208 10944 5234 10947
rect 5208 10915 5234 10918
rect 4748 10808 4774 10811
rect 4748 10779 4774 10782
rect 5122 10505 5136 10915
rect 5116 10502 5142 10505
rect 5116 10473 5142 10476
rect 5214 10403 5228 10915
rect 5352 10675 5366 11017
rect 5536 11015 5550 11187
rect 5628 11015 5642 11255
rect 5530 11012 5556 11015
rect 5530 10983 5556 10986
rect 5622 11012 5648 11015
rect 5622 10983 5648 10986
rect 5346 10672 5372 10675
rect 5346 10643 5372 10646
rect 5628 10573 5642 10983
rect 5622 10570 5648 10573
rect 5622 10541 5648 10544
rect 5208 10400 5234 10403
rect 5208 10371 5234 10374
rect 5214 5628 5228 10371
rect 5628 8839 5642 10541
rect 5674 10471 5688 12037
rect 5904 11865 5918 12063
rect 5898 11862 5924 11865
rect 5898 11833 5924 11836
rect 5904 11559 5918 11833
rect 5950 11559 5964 12071
rect 5898 11556 5924 11559
rect 5898 11527 5924 11530
rect 5944 11556 5970 11559
rect 5944 11527 5970 11530
rect 5760 11352 5786 11355
rect 5760 11323 5786 11326
rect 5766 11015 5780 11323
rect 5904 11287 5918 11527
rect 6134 11525 6148 14757
rect 6410 14075 6424 14995
rect 6456 14925 6470 15097
rect 6450 14922 6476 14925
rect 6450 14893 6476 14896
rect 6817 14600 6845 14604
rect 6817 14567 6818 14572
rect 6844 14567 6845 14572
rect 6818 14553 6844 14556
rect 6864 14480 6890 14483
rect 6864 14451 6890 14454
rect 6404 14072 6430 14075
rect 6404 14043 6430 14046
rect 6266 14038 6292 14041
rect 6266 14009 6292 14012
rect 6450 14038 6476 14041
rect 6450 14009 6476 14012
rect 6272 13837 6286 14009
rect 6312 13970 6338 13973
rect 6312 13941 6338 13944
rect 6266 13834 6292 13837
rect 6266 13805 6292 13808
rect 6318 13497 6332 13941
rect 6404 13936 6430 13939
rect 6404 13907 6430 13910
rect 6312 13494 6338 13497
rect 6312 13465 6338 13468
rect 6174 13392 6200 13395
rect 6174 13363 6200 13366
rect 6180 12953 6194 13363
rect 6318 12987 6332 13465
rect 6358 13120 6384 13123
rect 6358 13091 6384 13094
rect 6364 12987 6378 13091
rect 6312 12984 6338 12987
rect 6312 12955 6338 12958
rect 6358 12984 6384 12987
rect 6358 12955 6384 12958
rect 6174 12950 6200 12953
rect 6174 12921 6200 12924
rect 6220 12950 6246 12953
rect 6220 12921 6246 12924
rect 6226 12749 6240 12921
rect 6220 12746 6246 12749
rect 6220 12717 6246 12720
rect 6174 11556 6200 11559
rect 6174 11527 6200 11530
rect 6128 11522 6154 11525
rect 6128 11493 6154 11496
rect 6180 11355 6194 11527
rect 6174 11352 6200 11355
rect 6174 11323 6200 11326
rect 6410 11321 6424 13907
rect 6456 12987 6470 14009
rect 6870 13463 6884 14451
rect 6916 14381 6930 15097
rect 6910 14378 6936 14381
rect 6910 14349 6936 14352
rect 6962 14279 6976 15863
rect 7002 15330 7028 15333
rect 7002 15301 7028 15304
rect 7008 14823 7022 15301
rect 7054 15163 7068 16967
rect 7100 15333 7114 18361
rect 7284 18291 7298 18905
rect 7514 18333 7528 18939
rect 7468 18319 7528 18333
rect 7278 18288 7304 18291
rect 7278 18259 7304 18262
rect 7468 17339 7482 18319
rect 7508 18288 7534 18291
rect 7508 18259 7534 18262
rect 7514 18087 7528 18259
rect 7560 18121 7574 19483
rect 7554 18118 7580 18121
rect 7554 18089 7580 18092
rect 7652 18087 7666 20469
rect 7508 18084 7534 18087
rect 7508 18055 7534 18058
rect 7646 18084 7672 18087
rect 7646 18055 7672 18058
rect 7600 18050 7626 18053
rect 7600 18021 7626 18024
rect 7606 17815 7620 18021
rect 7600 17812 7626 17815
rect 7600 17783 7626 17786
rect 7652 17721 7666 18055
rect 7698 18019 7712 20469
rect 7790 20025 7804 20537
rect 7784 20022 7810 20025
rect 7784 19993 7810 19996
rect 7692 18016 7718 18019
rect 7692 17987 7718 17990
rect 7606 17707 7666 17721
rect 7462 17336 7488 17339
rect 7462 17307 7488 17310
rect 7232 17302 7258 17305
rect 7232 17273 7258 17276
rect 7140 16962 7166 16965
rect 7140 16933 7166 16936
rect 7094 15330 7120 15333
rect 7094 15301 7120 15304
rect 7146 15273 7160 16933
rect 7238 16455 7252 17273
rect 7468 16965 7482 17307
rect 7554 17302 7580 17305
rect 7554 17273 7580 17276
rect 7462 16962 7488 16965
rect 7462 16933 7488 16936
rect 7560 16761 7574 17273
rect 7554 16758 7580 16761
rect 7554 16729 7580 16732
rect 7278 16724 7304 16727
rect 7278 16695 7304 16698
rect 7284 16489 7298 16695
rect 7278 16486 7304 16489
rect 7278 16457 7304 16460
rect 7232 16452 7258 16455
rect 7232 16423 7258 16426
rect 7186 16418 7212 16421
rect 7186 16389 7212 16392
rect 7192 16149 7206 16389
rect 7284 16217 7298 16457
rect 7416 16452 7442 16455
rect 7416 16423 7442 16426
rect 7278 16214 7304 16217
rect 7278 16185 7304 16188
rect 7186 16146 7212 16149
rect 7186 16117 7212 16120
rect 7232 15840 7258 15843
rect 7232 15811 7258 15814
rect 7100 15259 7160 15273
rect 7048 15160 7074 15163
rect 7048 15131 7074 15134
rect 7002 14820 7028 14823
rect 7002 14791 7028 14794
rect 7100 14585 7114 15259
rect 7140 15194 7166 15197
rect 7140 15165 7166 15168
rect 7146 15148 7160 15165
rect 7139 15144 7167 15148
rect 7139 15111 7167 15116
rect 7094 14582 7120 14585
rect 7094 14553 7120 14556
rect 6956 14276 6982 14279
rect 6956 14247 6982 14250
rect 6956 13528 6982 13531
rect 6956 13499 6982 13502
rect 7186 13528 7212 13531
rect 7186 13499 7212 13502
rect 6864 13460 6890 13463
rect 6864 13431 6890 13434
rect 6450 12984 6476 12987
rect 6450 12955 6476 12958
rect 6496 12916 6522 12919
rect 6496 12887 6522 12890
rect 6502 12647 6516 12887
rect 6870 12851 6884 13431
rect 6962 12944 6976 13499
rect 7192 13312 7206 13499
rect 7185 13308 7213 13312
rect 7185 13275 7213 13280
rect 7094 12950 7120 12953
rect 6962 12930 7094 12944
rect 7094 12921 7120 12924
rect 6864 12848 6890 12851
rect 6864 12819 6890 12822
rect 6870 12681 6884 12819
rect 6864 12678 6890 12681
rect 6864 12649 6890 12652
rect 6496 12644 6522 12647
rect 6496 12615 6522 12618
rect 6542 12576 6568 12579
rect 6542 12547 6568 12550
rect 6548 12409 6562 12547
rect 6870 12409 6884 12649
rect 6909 12492 6937 12496
rect 6909 12459 6937 12464
rect 6916 12443 6930 12459
rect 6910 12440 6936 12443
rect 6910 12411 6936 12414
rect 6542 12406 6568 12409
rect 6542 12377 6568 12380
rect 6864 12406 6890 12409
rect 6864 12377 6890 12380
rect 6870 11831 6884 12377
rect 6864 11828 6890 11831
rect 6864 11799 6890 11802
rect 6863 11472 6891 11476
rect 6863 11439 6891 11444
rect 6870 11355 6884 11439
rect 6864 11352 6890 11355
rect 6864 11323 6890 11326
rect 6404 11318 6430 11321
rect 6404 11289 6430 11292
rect 5898 11284 5924 11287
rect 5898 11255 5924 11258
rect 6916 11015 6930 12411
rect 7100 12400 7114 12921
rect 7238 12647 7252 15811
rect 7422 15367 7436 16423
rect 7560 16225 7574 16729
rect 7514 16217 7574 16225
rect 7508 16214 7574 16217
rect 7534 16211 7574 16214
rect 7508 16185 7534 16188
rect 7514 15911 7528 16185
rect 7508 15908 7534 15911
rect 7508 15879 7534 15882
rect 7278 15364 7304 15367
rect 7278 15335 7304 15338
rect 7416 15364 7442 15367
rect 7416 15335 7442 15338
rect 7284 15095 7298 15335
rect 7606 15148 7620 17707
rect 7599 15144 7627 15148
rect 7324 15126 7350 15129
rect 7599 15111 7627 15116
rect 7324 15097 7350 15100
rect 7278 15092 7304 15095
rect 7278 15063 7304 15066
rect 7330 15069 7344 15097
rect 7284 14483 7298 15063
rect 7330 15055 7482 15069
rect 7468 15027 7482 15055
rect 7416 15024 7442 15027
rect 7416 14995 7442 14998
rect 7462 15024 7488 15027
rect 7462 14995 7488 14998
rect 7422 14823 7436 14995
rect 7698 14823 7712 17987
rect 7882 17305 7896 23691
rect 7928 21113 7942 24439
rect 8014 24413 8040 24416
rect 8066 24411 8080 24515
rect 8060 24408 8086 24411
rect 8060 24379 8086 24382
rect 7968 21280 7994 21283
rect 7968 21251 7994 21254
rect 7974 21113 7988 21251
rect 7922 21110 7948 21113
rect 7922 21081 7948 21084
rect 7968 21110 7994 21113
rect 7968 21081 7994 21084
rect 7922 21008 7948 21011
rect 7922 20979 7948 20982
rect 7928 20637 7942 20979
rect 7922 20634 7948 20637
rect 7922 20605 7948 20608
rect 7876 17302 7902 17305
rect 7876 17273 7902 17276
rect 8112 15367 8126 25603
rect 8526 25533 8540 25671
rect 8848 25533 8862 25943
rect 8520 25530 8546 25533
rect 8520 25501 8546 25504
rect 8658 25530 8684 25533
rect 8658 25501 8684 25504
rect 8842 25530 8868 25533
rect 8842 25501 8868 25504
rect 8336 25428 8362 25431
rect 8336 25399 8362 25402
rect 8152 25394 8178 25397
rect 8152 25365 8178 25368
rect 8158 25261 8172 25365
rect 8152 25258 8178 25261
rect 8152 25229 8178 25232
rect 8290 25156 8316 25159
rect 8290 25127 8316 25130
rect 8296 24912 8310 25127
rect 8342 25125 8356 25399
rect 8664 25159 8678 25501
rect 8940 25473 8954 26147
rect 9078 26043 9092 26419
rect 9072 26040 9098 26043
rect 9072 26011 9098 26014
rect 9124 25703 9138 28153
rect 9354 27335 9368 28663
rect 10228 28423 10242 29199
rect 10366 29069 10380 29479
rect 10360 29066 10386 29069
rect 10360 29037 10386 29040
rect 10406 28998 10432 29001
rect 10406 28969 10432 28972
rect 10360 28930 10386 28933
rect 10360 28901 10386 28904
rect 10366 28729 10380 28901
rect 10360 28726 10386 28729
rect 10360 28697 10386 28700
rect 10360 28624 10386 28627
rect 10360 28595 10386 28598
rect 10222 28420 10248 28423
rect 10222 28391 10248 28394
rect 10130 28386 10156 28389
rect 10130 28357 10156 28360
rect 10136 28117 10150 28357
rect 10176 28182 10202 28185
rect 10176 28153 10202 28156
rect 10130 28114 10156 28117
rect 10130 28085 10156 28088
rect 10182 27981 10196 28153
rect 10176 27978 10202 27981
rect 10176 27949 10202 27952
rect 9348 27332 9374 27335
rect 9348 27303 9374 27306
rect 9716 27332 9742 27335
rect 9716 27303 9742 27306
rect 9354 27131 9368 27303
rect 9348 27128 9374 27131
rect 9348 27099 9374 27102
rect 9722 27029 9736 27303
rect 9716 27026 9742 27029
rect 9716 26997 9742 27000
rect 9348 26992 9374 26995
rect 9348 26963 9374 26966
rect 9256 26550 9282 26553
rect 9256 26521 9282 26524
rect 9262 25907 9276 26521
rect 9354 26519 9368 26963
rect 10228 26791 10242 28391
rect 10366 28185 10380 28595
rect 10360 28182 10386 28185
rect 10360 28153 10386 28156
rect 10412 27879 10426 28969
rect 10504 28967 10518 29479
rect 10544 29440 10570 29443
rect 10544 29411 10570 29414
rect 10550 29171 10564 29411
rect 10544 29168 10570 29171
rect 10544 29139 10570 29142
rect 10550 29001 10564 29139
rect 11378 29069 11392 29479
rect 11878 29474 11904 29477
rect 11878 29445 11904 29448
rect 11648 29168 11674 29171
rect 11648 29139 11674 29142
rect 11372 29066 11398 29069
rect 11372 29037 11398 29040
rect 10544 28998 10570 29001
rect 10544 28969 10570 28972
rect 10498 28964 10524 28967
rect 10498 28935 10524 28938
rect 10504 28763 10518 28935
rect 10550 28933 10564 28969
rect 11654 28967 11668 29139
rect 11884 29069 11898 29445
rect 12108 29440 12134 29443
rect 12108 29411 12134 29414
rect 12114 29307 12128 29411
rect 12108 29304 12134 29307
rect 12108 29275 12134 29278
rect 11878 29066 11904 29069
rect 11878 29037 11904 29040
rect 11188 28964 11214 28967
rect 11188 28935 11214 28938
rect 11648 28964 11674 28967
rect 11648 28935 11674 28938
rect 11786 28964 11812 28967
rect 11786 28935 11812 28938
rect 10544 28930 10570 28933
rect 10544 28901 10570 28904
rect 10498 28760 10524 28763
rect 10498 28731 10524 28734
rect 10504 28185 10518 28731
rect 10550 28253 10564 28901
rect 11194 28729 11208 28935
rect 11188 28726 11214 28729
rect 11188 28697 11214 28700
rect 10866 28352 10892 28355
rect 10866 28323 10892 28326
rect 10544 28250 10570 28253
rect 10544 28221 10570 28224
rect 10498 28182 10524 28185
rect 10498 28153 10524 28156
rect 10872 28151 10886 28323
rect 11194 28253 11208 28697
rect 11188 28250 11214 28253
rect 11188 28221 11214 28224
rect 11792 28219 11806 28935
rect 11786 28216 11812 28219
rect 11786 28187 11812 28190
rect 12246 28216 12272 28219
rect 12246 28187 12272 28190
rect 11004 28182 11030 28185
rect 11004 28153 11030 28156
rect 10866 28148 10892 28151
rect 10866 28119 10892 28122
rect 10498 28080 10524 28083
rect 10498 28051 10524 28054
rect 10504 27879 10518 28051
rect 10406 27876 10432 27879
rect 10406 27847 10432 27850
rect 10498 27876 10524 27879
rect 10498 27847 10524 27850
rect 10268 27638 10294 27641
rect 10268 27609 10294 27612
rect 10274 27369 10288 27609
rect 10412 27573 10426 27847
rect 10406 27570 10432 27573
rect 10406 27541 10432 27544
rect 10268 27366 10294 27369
rect 10268 27337 10294 27340
rect 10222 26788 10248 26791
rect 10222 26759 10248 26762
rect 10504 26519 10518 27847
rect 10544 27672 10570 27675
rect 10544 27643 10570 27646
rect 10550 26723 10564 27643
rect 11010 27641 11024 28153
rect 11694 28148 11720 28151
rect 11694 28119 11720 28122
rect 11648 27876 11674 27879
rect 11648 27847 11674 27850
rect 11602 27808 11628 27811
rect 11602 27779 11628 27782
rect 11004 27638 11030 27641
rect 11004 27609 11030 27612
rect 10636 27570 10662 27573
rect 10636 27541 10662 27544
rect 10642 27131 10656 27541
rect 10636 27128 10662 27131
rect 10636 27099 10662 27102
rect 10728 27128 10754 27131
rect 10728 27099 10754 27102
rect 10544 26720 10570 26723
rect 10544 26691 10570 26694
rect 10550 26553 10564 26691
rect 10734 26621 10748 27099
rect 11608 27029 11622 27779
rect 11654 27675 11668 27847
rect 11648 27672 11674 27675
rect 11648 27643 11674 27646
rect 11700 27641 11714 28119
rect 11792 27879 11806 28187
rect 11786 27876 11812 27879
rect 11786 27847 11812 27850
rect 12108 27876 12134 27879
rect 12108 27847 12134 27850
rect 12114 27709 12128 27847
rect 12108 27706 12134 27709
rect 12108 27677 12134 27680
rect 12114 27641 12128 27677
rect 12252 27641 12266 28187
rect 11694 27638 11720 27641
rect 11694 27609 11720 27612
rect 11924 27638 11950 27641
rect 11924 27609 11950 27612
rect 12108 27638 12134 27641
rect 12108 27609 12134 27612
rect 12246 27638 12272 27641
rect 12246 27609 12272 27612
rect 11930 27165 11944 27609
rect 11924 27162 11950 27165
rect 11924 27133 11950 27136
rect 12298 27097 12312 29479
rect 12338 29474 12364 29477
rect 12338 29445 12364 29448
rect 12344 27607 12358 29445
rect 13810 29270 13836 29273
rect 13810 29241 13836 29244
rect 13120 29236 13146 29239
rect 13120 29207 13146 29210
rect 13126 29035 13140 29207
rect 13816 29069 13830 29241
rect 13948 29202 13974 29205
rect 13948 29173 13974 29176
rect 13902 29168 13928 29171
rect 13902 29139 13928 29142
rect 13810 29066 13836 29069
rect 13810 29037 13836 29040
rect 13120 29032 13146 29035
rect 13120 29003 13146 29006
rect 13074 28386 13100 28389
rect 13074 28357 13100 28360
rect 13080 28253 13094 28357
rect 13126 28355 13140 29003
rect 13908 29001 13922 29139
rect 13902 28998 13928 29001
rect 13902 28969 13928 28972
rect 13258 28692 13284 28695
rect 13258 28663 13284 28666
rect 13212 28658 13238 28661
rect 13212 28629 13238 28632
rect 13218 28389 13232 28629
rect 13212 28386 13238 28389
rect 13212 28357 13238 28360
rect 13120 28352 13146 28355
rect 13120 28323 13146 28326
rect 13074 28250 13100 28253
rect 13074 28221 13100 28224
rect 12384 28182 12410 28185
rect 12384 28153 12410 28156
rect 12390 27879 12404 28153
rect 12384 27876 12410 27879
rect 12384 27847 12410 27850
rect 12338 27604 12364 27607
rect 12338 27575 12364 27578
rect 12390 27131 12404 27847
rect 13126 27335 13140 28323
rect 13264 27607 13278 28663
rect 13304 28624 13330 28627
rect 13304 28595 13330 28598
rect 13310 28185 13324 28595
rect 13304 28182 13330 28185
rect 13304 28153 13330 28156
rect 13350 27638 13376 27641
rect 13350 27609 13376 27612
rect 13396 27638 13422 27641
rect 13396 27609 13422 27612
rect 13580 27638 13606 27641
rect 13580 27609 13606 27612
rect 13264 27593 13324 27607
rect 13310 27573 13324 27593
rect 13304 27570 13330 27573
rect 13304 27541 13330 27544
rect 13258 27536 13284 27539
rect 13258 27507 13284 27510
rect 13264 27335 13278 27507
rect 13120 27332 13146 27335
rect 13120 27303 13146 27306
rect 13258 27332 13284 27335
rect 13258 27303 13284 27306
rect 12384 27128 12410 27131
rect 12384 27099 12410 27102
rect 11924 27094 11950 27097
rect 11924 27065 11950 27068
rect 12292 27094 12318 27097
rect 12292 27065 12318 27068
rect 11930 27037 11944 27065
rect 11602 27026 11628 27029
rect 11930 27023 11990 27037
rect 11602 26997 11628 27000
rect 10820 26992 10846 26995
rect 10820 26963 10846 26966
rect 10826 26791 10840 26963
rect 10820 26788 10846 26791
rect 10820 26759 10846 26762
rect 11050 26754 11076 26757
rect 11050 26725 11076 26728
rect 10728 26618 10754 26621
rect 10728 26589 10754 26592
rect 10544 26550 10570 26553
rect 10544 26521 10570 26524
rect 9302 26516 9328 26519
rect 9302 26487 9328 26490
rect 9348 26516 9374 26519
rect 9348 26487 9374 26490
rect 10498 26516 10524 26519
rect 10498 26487 10524 26490
rect 9308 26281 9322 26487
rect 10820 26312 10846 26315
rect 10820 26283 10846 26286
rect 9302 26278 9328 26281
rect 9302 26249 9328 26252
rect 9256 25904 9282 25907
rect 9256 25875 9282 25878
rect 10130 25904 10156 25907
rect 10130 25875 10156 25878
rect 9262 25805 9276 25875
rect 9256 25802 9282 25805
rect 9256 25773 9282 25776
rect 9118 25700 9144 25703
rect 9118 25671 9144 25674
rect 9578 25700 9604 25703
rect 9578 25671 9604 25674
rect 8940 25465 9092 25473
rect 8940 25462 9098 25465
rect 8940 25459 9072 25462
rect 8940 25431 8954 25459
rect 9072 25433 9098 25436
rect 8934 25428 8960 25431
rect 8934 25399 8960 25402
rect 8658 25156 8684 25159
rect 8658 25127 8684 25130
rect 8336 25122 8362 25125
rect 8336 25093 8362 25096
rect 8204 24898 8310 24912
rect 8204 24615 8218 24898
rect 8198 24612 8224 24615
rect 8244 24612 8270 24615
rect 8198 24583 8224 24586
rect 8243 24596 8244 24600
rect 8270 24596 8271 24600
rect 8204 24173 8218 24583
rect 8243 24563 8271 24568
rect 8244 24544 8270 24547
rect 8342 24521 8356 25093
rect 8940 24921 8954 25399
rect 8934 24918 8960 24921
rect 8934 24889 8960 24892
rect 9210 24612 9236 24615
rect 9210 24583 9236 24586
rect 8270 24518 8356 24521
rect 8244 24515 8356 24518
rect 8250 24507 8356 24515
rect 8198 24170 8224 24173
rect 8198 24141 8224 24144
rect 8204 23569 8218 24141
rect 8342 24071 8356 24507
rect 9164 24374 9190 24377
rect 9164 24345 9190 24348
rect 9170 24173 9184 24345
rect 9216 24173 9230 24583
rect 9302 24544 9328 24547
rect 9302 24515 9328 24518
rect 9308 24411 9322 24515
rect 9302 24408 9328 24411
rect 9302 24379 9328 24382
rect 9256 24374 9282 24377
rect 9256 24345 9282 24348
rect 9348 24374 9374 24377
rect 9348 24345 9374 24348
rect 9164 24170 9190 24173
rect 9164 24141 9190 24144
rect 9210 24170 9236 24173
rect 9210 24141 9236 24144
rect 9262 24157 9276 24345
rect 9354 24275 9368 24345
rect 9440 24340 9466 24343
rect 9440 24311 9466 24314
rect 9348 24272 9374 24275
rect 9348 24243 9374 24246
rect 9262 24143 9322 24157
rect 9026 24136 9052 24139
rect 9026 24107 9052 24110
rect 8336 24068 8362 24071
rect 8336 24039 8362 24042
rect 8381 24052 8409 24056
rect 8342 23569 8356 24039
rect 8381 24019 8409 24024
rect 8158 23555 8218 23569
rect 8296 23555 8356 23569
rect 8158 23527 8172 23555
rect 8296 23527 8310 23555
rect 8152 23524 8178 23527
rect 8152 23495 8178 23498
rect 8290 23524 8316 23527
rect 8290 23495 8316 23498
rect 8388 23493 8402 24019
rect 9032 23833 9046 24107
rect 9164 24068 9190 24071
rect 9164 24039 9190 24042
rect 9170 23833 9184 24039
rect 9026 23830 9052 23833
rect 9026 23801 9052 23804
rect 9164 23830 9190 23833
rect 9164 23801 9190 23804
rect 8888 23524 8914 23527
rect 8887 23508 8888 23512
rect 8914 23508 8915 23512
rect 8382 23490 8408 23493
rect 8887 23475 8915 23480
rect 8382 23461 8408 23464
rect 8198 23456 8224 23459
rect 8224 23430 8310 23433
rect 8198 23427 8310 23430
rect 8204 23419 8310 23427
rect 8296 22541 8310 23419
rect 8658 22640 8684 22643
rect 8658 22611 8684 22614
rect 8290 22538 8316 22541
rect 8290 22509 8316 22512
rect 8664 22507 8678 22611
rect 8658 22504 8684 22507
rect 8658 22475 8684 22478
rect 8336 22470 8362 22473
rect 8336 22441 8362 22444
rect 8290 21552 8316 21555
rect 8290 21523 8316 21526
rect 8296 21419 8310 21523
rect 8290 21416 8316 21419
rect 8290 21387 8316 21390
rect 8244 21348 8270 21351
rect 8244 21319 8270 21322
rect 8250 21172 8264 21319
rect 8342 21283 8356 22441
rect 8428 22402 8454 22405
rect 8428 22373 8454 22376
rect 8434 22269 8448 22373
rect 8428 22266 8454 22269
rect 8428 22237 8454 22240
rect 8520 21688 8546 21691
rect 8520 21659 8546 21662
rect 8526 21453 8540 21659
rect 8520 21450 8546 21453
rect 8520 21421 8546 21424
rect 8336 21280 8362 21283
rect 8336 21251 8362 21254
rect 8290 21178 8316 21181
rect 8250 21158 8290 21172
rect 8290 21149 8316 21152
rect 8342 20707 8356 21251
rect 8342 20693 8402 20707
rect 8290 20566 8316 20569
rect 8290 20537 8316 20540
rect 8244 19410 8270 19413
rect 8244 19381 8270 19384
rect 8250 19277 8264 19381
rect 8244 19274 8270 19277
rect 8244 19245 8270 19248
rect 8296 19175 8310 20537
rect 8388 19481 8402 20693
rect 8382 19478 8408 19481
rect 8382 19449 8408 19452
rect 8290 19172 8316 19175
rect 8290 19143 8316 19146
rect 8474 19172 8500 19175
rect 8474 19143 8500 19146
rect 8290 18628 8316 18631
rect 8290 18599 8316 18602
rect 8296 18087 8310 18599
rect 8290 18084 8316 18087
rect 8290 18055 8316 18058
rect 8428 18084 8454 18087
rect 8428 18055 8454 18058
rect 8336 18050 8362 18053
rect 8336 18021 8362 18024
rect 8290 17200 8316 17203
rect 8290 17171 8316 17174
rect 8244 16214 8270 16217
rect 8244 16185 8270 16188
rect 8198 16112 8224 16115
rect 8198 16083 8224 16086
rect 8204 15911 8218 16083
rect 8198 15908 8224 15911
rect 8198 15879 8224 15882
rect 8250 15885 8264 16185
rect 8296 15979 8310 17171
rect 8342 16761 8356 18021
rect 8434 17645 8448 18055
rect 8428 17642 8454 17645
rect 8428 17613 8454 17616
rect 8434 17237 8448 17613
rect 8480 17509 8494 19143
rect 8526 18597 8540 21421
rect 8658 21348 8684 21351
rect 8658 21319 8684 21322
rect 8612 21280 8638 21283
rect 8612 21251 8638 21254
rect 8618 20909 8632 21251
rect 8664 21079 8678 21319
rect 8894 21317 8908 23475
rect 9032 23255 9046 23801
rect 9170 23289 9184 23801
rect 9164 23286 9190 23289
rect 9164 23257 9190 23260
rect 9026 23252 9052 23255
rect 9026 23223 9052 23226
rect 9032 22711 9046 23223
rect 9026 22708 9052 22711
rect 9026 22679 9052 22682
rect 8980 22368 9006 22371
rect 8980 22339 9006 22342
rect 8888 21314 8914 21317
rect 8888 21285 8914 21288
rect 8704 21280 8730 21283
rect 8704 21251 8730 21254
rect 8710 21113 8724 21251
rect 8704 21110 8730 21113
rect 8704 21081 8730 21084
rect 8658 21076 8684 21079
rect 8658 21047 8684 21050
rect 8612 20906 8638 20909
rect 8612 20877 8638 20880
rect 8664 20025 8678 21047
rect 8986 20501 9000 22339
rect 9032 22201 9046 22679
rect 9072 22436 9098 22439
rect 9072 22407 9098 22410
rect 9026 22198 9052 22201
rect 9026 22169 9052 22172
rect 9078 21351 9092 22407
rect 9216 22277 9230 24141
rect 9256 23320 9282 23323
rect 9256 23291 9282 23294
rect 9262 23017 9276 23291
rect 9256 23014 9282 23017
rect 9256 22985 9282 22988
rect 9262 22915 9276 22985
rect 9256 22912 9282 22915
rect 9256 22883 9282 22886
rect 9170 22263 9230 22277
rect 9170 22235 9184 22263
rect 9164 22232 9190 22235
rect 9164 22203 9190 22206
rect 9308 21453 9322 24143
rect 9446 23527 9460 24311
rect 9440 23524 9466 23527
rect 9440 23495 9466 23498
rect 9532 23524 9558 23527
rect 9532 23495 9558 23498
rect 9394 23456 9420 23459
rect 9394 23427 9420 23430
rect 9348 23286 9374 23289
rect 9348 23257 9374 23260
rect 9354 22745 9368 23257
rect 9400 22983 9414 23427
rect 9538 23085 9552 23495
rect 9532 23082 9558 23085
rect 9532 23053 9558 23056
rect 9394 22980 9420 22983
rect 9394 22951 9420 22954
rect 9348 22742 9374 22745
rect 9348 22713 9374 22716
rect 9302 21450 9328 21453
rect 9302 21421 9328 21424
rect 9072 21348 9098 21351
rect 9072 21319 9098 21322
rect 9078 20707 9092 21319
rect 9078 20693 9138 20707
rect 8980 20498 9006 20501
rect 8980 20469 9006 20472
rect 9026 20362 9052 20365
rect 9026 20333 9052 20336
rect 9032 20195 9046 20333
rect 9026 20192 9052 20195
rect 9026 20163 9052 20166
rect 9032 20059 9046 20163
rect 9026 20056 9052 20059
rect 9026 20027 9052 20030
rect 8658 20022 8684 20025
rect 8658 19993 8684 19996
rect 9072 20022 9098 20025
rect 9072 19993 9098 19996
rect 8664 19753 8678 19993
rect 8658 19750 8684 19753
rect 8658 19721 8684 19724
rect 9078 19719 9092 19993
rect 9072 19716 9098 19719
rect 8703 19700 8731 19704
rect 9072 19687 9098 19690
rect 8703 19667 8704 19672
rect 8730 19667 8731 19672
rect 8704 19653 8730 19656
rect 8842 19478 8868 19481
rect 8842 19449 8868 19452
rect 8848 19277 8862 19449
rect 8980 19410 9006 19413
rect 8980 19381 9006 19384
rect 8842 19274 8868 19277
rect 8842 19245 8868 19248
rect 8986 19005 9000 19381
rect 8980 19002 9006 19005
rect 8980 18973 9006 18976
rect 9078 18835 9092 19687
rect 9124 19481 9138 20693
rect 9308 19914 9322 21421
rect 9354 20025 9368 22713
rect 9584 20909 9598 25671
rect 9624 25530 9650 25533
rect 9624 25501 9650 25504
rect 9630 25363 9644 25501
rect 9624 25360 9650 25363
rect 9624 25331 9650 25334
rect 9630 24887 9644 25331
rect 9670 24952 9696 24955
rect 9670 24923 9696 24926
rect 9624 24884 9650 24887
rect 9624 24855 9650 24858
rect 9624 24272 9650 24275
rect 9624 24243 9650 24246
rect 9630 22269 9644 24243
rect 9676 23988 9690 24923
rect 9669 23984 9697 23988
rect 9669 23951 9697 23956
rect 9676 23731 9690 23951
rect 9670 23728 9696 23731
rect 9670 23699 9696 23702
rect 9716 22776 9742 22779
rect 9716 22747 9742 22750
rect 9670 22708 9696 22711
rect 9670 22679 9696 22682
rect 9624 22266 9650 22269
rect 9624 22237 9650 22240
rect 9676 21657 9690 22679
rect 9722 21997 9736 22747
rect 9808 22198 9834 22201
rect 9808 22169 9834 22172
rect 9716 21994 9742 21997
rect 9716 21965 9742 21968
rect 9670 21654 9696 21657
rect 9670 21625 9696 21628
rect 9676 21283 9690 21625
rect 9670 21280 9696 21283
rect 9670 21251 9696 21254
rect 9676 21011 9690 21251
rect 9722 21138 9736 21965
rect 9814 21657 9828 22169
rect 9899 21808 9927 21812
rect 9899 21775 9927 21780
rect 9906 21691 9920 21775
rect 9900 21688 9926 21691
rect 9900 21659 9926 21662
rect 9808 21654 9834 21657
rect 9808 21625 9834 21628
rect 9762 21144 9788 21147
rect 9722 21124 9762 21138
rect 9762 21115 9788 21118
rect 9814 21113 9828 21625
rect 9808 21110 9834 21113
rect 9808 21081 9834 21084
rect 9670 21008 9696 21011
rect 9670 20979 9696 20982
rect 9578 20906 9604 20909
rect 9578 20877 9604 20880
rect 9348 20022 9374 20025
rect 9348 19993 9374 19996
rect 10084 20022 10110 20025
rect 10084 19993 10110 19996
rect 9348 19920 9374 19923
rect 9308 19900 9348 19914
rect 9118 19478 9144 19481
rect 9118 19449 9144 19452
rect 9210 19478 9236 19481
rect 9210 19449 9236 19452
rect 8566 18832 8592 18835
rect 8566 18803 8592 18806
rect 9072 18832 9098 18835
rect 9072 18803 9098 18806
rect 8572 18631 8586 18803
rect 8566 18628 8592 18631
rect 8566 18599 8592 18602
rect 8520 18594 8546 18597
rect 8520 18565 8546 18568
rect 8572 18087 8586 18599
rect 9216 18291 9230 19449
rect 9308 19447 9322 19900
rect 9348 19891 9374 19894
rect 10090 19821 10104 19993
rect 10084 19818 10110 19821
rect 10084 19789 10110 19792
rect 9578 19750 9604 19753
rect 9578 19721 9604 19724
rect 9302 19444 9328 19447
rect 9302 19415 9328 19418
rect 9302 19376 9328 19379
rect 9302 19347 9328 19350
rect 9308 18393 9322 19347
rect 9584 19327 9598 19721
rect 9624 19444 9650 19447
rect 9624 19415 9650 19418
rect 9446 19313 9598 19327
rect 9348 18628 9374 18631
rect 9348 18599 9374 18602
rect 9302 18390 9328 18393
rect 9302 18361 9328 18364
rect 9210 18288 9236 18291
rect 9210 18259 9236 18262
rect 9118 18186 9144 18189
rect 9144 18166 9184 18180
rect 9118 18157 9144 18160
rect 8566 18084 8592 18087
rect 8566 18055 8592 18058
rect 8572 17543 8586 18055
rect 8566 17540 8592 17543
rect 8566 17511 8592 17514
rect 8474 17506 8500 17509
rect 8474 17477 8500 17480
rect 8428 17234 8454 17237
rect 8428 17205 8454 17208
rect 8336 16758 8362 16761
rect 8336 16729 8362 16732
rect 8428 16758 8454 16761
rect 8428 16729 8454 16732
rect 8382 16724 8408 16727
rect 8342 16698 8382 16701
rect 8342 16695 8408 16698
rect 8342 16687 8402 16695
rect 8290 15976 8316 15979
rect 8290 15947 8316 15950
rect 8250 15871 8310 15885
rect 8244 15840 8270 15843
rect 8244 15811 8270 15814
rect 8106 15364 8132 15367
rect 8106 15335 8132 15338
rect 7784 15330 7810 15333
rect 7784 15301 7810 15304
rect 7790 15120 7804 15301
rect 7830 15126 7856 15129
rect 7790 15106 7830 15120
rect 7416 14820 7442 14823
rect 7416 14791 7442 14794
rect 7462 14820 7488 14823
rect 7462 14791 7488 14794
rect 7692 14820 7718 14823
rect 7692 14791 7718 14794
rect 7468 14653 7482 14791
rect 7462 14650 7488 14653
rect 7462 14621 7488 14624
rect 7790 14604 7804 15106
rect 7830 15097 7856 15100
rect 8250 14789 8264 15811
rect 8296 14823 8310 15871
rect 8342 15843 8356 16687
rect 8382 16656 8408 16659
rect 8382 16627 8408 16630
rect 8388 15843 8402 16627
rect 8336 15840 8362 15843
rect 8336 15811 8362 15814
rect 8382 15840 8408 15843
rect 8382 15811 8408 15814
rect 8434 15707 8448 16729
rect 8480 16217 8494 17477
rect 8658 17234 8684 17237
rect 8658 17205 8684 17208
rect 8664 17033 8678 17205
rect 8658 17030 8684 17033
rect 8658 17001 8684 17004
rect 8664 16769 8678 17001
rect 8980 16996 9006 16999
rect 8980 16967 9006 16970
rect 8934 16962 8960 16965
rect 8934 16933 8960 16936
rect 8940 16795 8954 16933
rect 8618 16755 8678 16769
rect 8934 16792 8960 16795
rect 8934 16763 8960 16766
rect 8618 16455 8632 16755
rect 8612 16452 8638 16455
rect 8612 16423 8638 16426
rect 8618 16217 8632 16423
rect 8934 16418 8960 16421
rect 8986 16412 9000 16967
rect 8960 16398 9000 16412
rect 8934 16389 8960 16392
rect 8986 16225 9000 16398
rect 9025 16300 9053 16304
rect 9025 16267 9053 16272
rect 9032 16251 9046 16267
rect 8940 16217 9000 16225
rect 9026 16248 9052 16251
rect 9026 16219 9052 16222
rect 8474 16214 8500 16217
rect 8474 16185 8500 16188
rect 8612 16214 8638 16217
rect 8612 16185 8638 16188
rect 8934 16214 9000 16217
rect 8960 16211 9000 16214
rect 8934 16185 8960 16188
rect 8986 16157 9000 16211
rect 8986 16143 9046 16157
rect 8980 16010 9006 16013
rect 8980 15981 9006 15984
rect 8428 15704 8454 15707
rect 8428 15675 8454 15678
rect 8434 15367 8448 15675
rect 8428 15364 8454 15367
rect 8428 15335 8454 15338
rect 8986 15197 9000 15981
rect 9032 15673 9046 16143
rect 9026 15670 9052 15673
rect 9026 15641 9052 15644
rect 9118 15636 9144 15639
rect 9118 15607 9144 15610
rect 9072 15296 9098 15299
rect 9072 15267 9098 15270
rect 9078 15197 9092 15267
rect 8980 15194 9006 15197
rect 8980 15165 9006 15168
rect 9072 15194 9098 15197
rect 9072 15165 9098 15168
rect 8842 15126 8868 15129
rect 8842 15097 8868 15100
rect 8290 14820 8316 14823
rect 8290 14791 8316 14794
rect 8520 14820 8546 14823
rect 8520 14791 8546 14794
rect 8244 14786 8270 14789
rect 8244 14757 8270 14760
rect 7783 14600 7811 14604
rect 7783 14567 7811 14572
rect 7278 14480 7304 14483
rect 7278 14451 7304 14454
rect 7284 14313 7298 14451
rect 7278 14310 7304 14313
rect 7278 14281 7304 14284
rect 7646 14310 7672 14313
rect 7646 14281 7672 14284
rect 7652 13769 7666 14281
rect 7790 14279 7804 14567
rect 8526 14551 8540 14791
rect 8704 14786 8730 14789
rect 8704 14757 8730 14760
rect 8520 14548 8546 14551
rect 7921 14532 7949 14536
rect 8520 14519 8546 14522
rect 7921 14499 7949 14504
rect 7784 14276 7810 14279
rect 7784 14247 7810 14250
rect 7646 13766 7672 13769
rect 7646 13737 7672 13740
rect 7928 13191 7942 14499
rect 8526 14497 8540 14519
rect 8480 14483 8540 14497
rect 8480 13769 8494 14483
rect 8710 14279 8724 14757
rect 8848 14381 8862 15097
rect 8888 15058 8914 15061
rect 8888 15029 8914 15032
rect 8894 14789 8908 15029
rect 8986 14823 9000 15165
rect 9124 15027 9138 15607
rect 9170 15095 9184 18166
rect 9216 15911 9230 18259
rect 9308 16013 9322 18361
rect 9302 16010 9328 16013
rect 9302 15981 9328 15984
rect 9210 15908 9236 15911
rect 9210 15879 9236 15882
rect 9216 15129 9230 15879
rect 9354 15877 9368 18599
rect 9394 18390 9420 18393
rect 9394 18361 9420 18364
rect 9400 17645 9414 18361
rect 9446 18325 9460 19313
rect 9532 18832 9558 18835
rect 9532 18803 9558 18806
rect 9486 18560 9512 18563
rect 9486 18531 9512 18534
rect 9492 18393 9506 18531
rect 9538 18461 9552 18803
rect 9532 18458 9558 18461
rect 9532 18429 9558 18432
rect 9531 18408 9559 18412
rect 9559 18400 9573 18403
rect 9486 18390 9512 18393
rect 9531 18375 9547 18380
rect 9547 18371 9573 18374
rect 9486 18361 9512 18364
rect 9440 18322 9466 18325
rect 9440 18293 9466 18296
rect 9486 18322 9512 18325
rect 9486 18293 9512 18296
rect 9492 18189 9506 18293
rect 9486 18186 9512 18189
rect 9486 18157 9512 18160
rect 9394 17642 9420 17645
rect 9394 17613 9420 17616
rect 9630 17203 9644 19415
rect 10038 17234 10064 17237
rect 10038 17205 10064 17208
rect 9624 17200 9650 17203
rect 9624 17171 9650 17174
rect 9532 16928 9558 16931
rect 9532 16899 9558 16902
rect 9538 16761 9552 16899
rect 9630 16761 9644 17171
rect 10044 16761 10058 17205
rect 10136 16965 10150 25875
rect 10682 25462 10708 25465
rect 10682 25433 10708 25436
rect 10498 25088 10524 25091
rect 10498 25059 10524 25062
rect 10504 24615 10518 25059
rect 10688 24955 10702 25433
rect 10774 25360 10800 25363
rect 10774 25331 10800 25334
rect 10682 24952 10708 24955
rect 10682 24923 10708 24926
rect 10636 24816 10662 24819
rect 10636 24787 10662 24790
rect 10543 24664 10571 24668
rect 10543 24631 10571 24636
rect 10550 24615 10564 24631
rect 10642 24615 10656 24787
rect 10780 24683 10794 25331
rect 10728 24680 10754 24683
rect 10728 24651 10754 24654
rect 10774 24680 10800 24683
rect 10774 24651 10800 24654
rect 10498 24612 10524 24615
rect 10498 24583 10524 24586
rect 10544 24612 10570 24615
rect 10544 24583 10570 24586
rect 10636 24612 10662 24615
rect 10636 24583 10662 24586
rect 10550 24377 10564 24583
rect 10682 24544 10708 24547
rect 10682 24515 10708 24518
rect 10544 24374 10570 24377
rect 10544 24345 10570 24348
rect 10222 23728 10248 23731
rect 10222 23699 10248 23702
rect 10228 23527 10242 23699
rect 10222 23524 10248 23527
rect 10222 23495 10248 23498
rect 10406 23524 10432 23527
rect 10406 23495 10432 23498
rect 10360 23490 10386 23493
rect 10360 23461 10386 23464
rect 10366 23357 10380 23461
rect 10360 23354 10386 23357
rect 10360 23325 10386 23328
rect 10412 23323 10426 23495
rect 10636 23456 10662 23459
rect 10636 23427 10662 23430
rect 10406 23320 10432 23323
rect 10406 23291 10432 23294
rect 10412 23187 10426 23291
rect 10642 23289 10656 23427
rect 10688 23357 10702 24515
rect 10734 24445 10748 24651
rect 10728 24442 10754 24445
rect 10728 24413 10754 24416
rect 10826 23357 10840 26283
rect 11056 25397 11070 26725
rect 11608 26247 11622 26997
rect 11878 26992 11904 26995
rect 11878 26963 11904 26966
rect 11884 26791 11898 26963
rect 11878 26788 11904 26791
rect 11878 26759 11904 26762
rect 11740 26754 11766 26757
rect 11740 26725 11766 26728
rect 11746 26553 11760 26725
rect 11976 26723 11990 27023
rect 12298 26791 12312 27065
rect 12200 26788 12226 26791
rect 12200 26759 12226 26762
rect 12292 26788 12318 26791
rect 12292 26759 12318 26762
rect 11970 26720 11996 26723
rect 11970 26691 11996 26694
rect 11740 26550 11766 26553
rect 11740 26521 11766 26524
rect 11602 26244 11628 26247
rect 11602 26215 11628 26218
rect 11050 25394 11076 25397
rect 11050 25365 11076 25368
rect 11004 25156 11030 25159
rect 11056 25133 11070 25365
rect 11234 25258 11260 25261
rect 11234 25229 11260 25232
rect 11030 25130 11070 25133
rect 11004 25127 11070 25130
rect 11010 25119 11070 25127
rect 11240 25125 11254 25229
rect 11326 25156 11352 25159
rect 11352 25136 11392 25150
rect 11326 25127 11352 25130
rect 11056 24887 11070 25119
rect 11234 25122 11260 25125
rect 11234 25093 11260 25096
rect 11378 24921 11392 25136
rect 11372 24918 11398 24921
rect 11372 24889 11398 24892
rect 11050 24884 11076 24887
rect 11050 24855 11076 24858
rect 11056 24615 11070 24855
rect 11326 24816 11352 24819
rect 11326 24787 11352 24790
rect 11050 24612 11076 24615
rect 11050 24583 11076 24586
rect 10958 23762 10984 23765
rect 10958 23733 10984 23736
rect 10964 23561 10978 23733
rect 11056 23569 11070 24583
rect 11332 24581 11346 24787
rect 11378 24615 11392 24889
rect 11372 24612 11398 24615
rect 11372 24583 11398 24586
rect 11326 24578 11352 24581
rect 11326 24549 11352 24552
rect 11332 23833 11346 24549
rect 11326 23830 11352 23833
rect 11326 23801 11352 23804
rect 10958 23558 10984 23561
rect 10958 23529 10984 23532
rect 11010 23555 11070 23569
rect 11010 23527 11024 23555
rect 11004 23524 11030 23527
rect 11004 23495 11030 23498
rect 10682 23354 10708 23357
rect 10682 23325 10708 23328
rect 10728 23354 10754 23357
rect 10728 23325 10754 23328
rect 10820 23354 10846 23357
rect 10820 23325 10846 23328
rect 10636 23286 10662 23289
rect 10636 23257 10662 23260
rect 10406 23184 10432 23187
rect 10406 23155 10432 23158
rect 10268 22946 10294 22949
rect 10268 22917 10294 22920
rect 10274 22832 10288 22917
rect 10267 22828 10295 22832
rect 10267 22795 10295 22800
rect 10274 21895 10288 22795
rect 10360 22266 10386 22269
rect 10360 22237 10386 22240
rect 10314 22096 10340 22099
rect 10314 22067 10340 22070
rect 10320 21895 10334 22067
rect 10366 21948 10380 22237
rect 10359 21944 10387 21948
rect 10359 21911 10387 21916
rect 10366 21895 10380 21911
rect 10176 21892 10202 21895
rect 10176 21863 10202 21866
rect 10268 21892 10294 21895
rect 10268 21863 10294 21866
rect 10314 21892 10340 21895
rect 10314 21863 10340 21866
rect 10360 21892 10386 21895
rect 10360 21863 10386 21866
rect 10182 21453 10196 21863
rect 10590 21824 10616 21827
rect 10590 21795 10616 21798
rect 10176 21450 10202 21453
rect 10176 21421 10202 21424
rect 10596 21351 10610 21795
rect 10590 21348 10616 21351
rect 10590 21319 10616 21322
rect 10636 21348 10662 21351
rect 10636 21319 10662 21322
rect 10314 21280 10340 21283
rect 10314 21251 10340 21254
rect 10222 21008 10248 21011
rect 10222 20979 10248 20982
rect 10228 20792 10242 20979
rect 10320 20841 10334 21251
rect 10642 21181 10656 21319
rect 10636 21178 10662 21181
rect 10636 21149 10662 21152
rect 10314 20838 10340 20841
rect 10314 20809 10340 20812
rect 10221 20788 10249 20792
rect 10221 20755 10249 20760
rect 10176 20498 10202 20501
rect 10176 20469 10202 20472
rect 10182 20059 10196 20469
rect 10176 20056 10202 20059
rect 10176 20027 10202 20030
rect 10228 18427 10242 20755
rect 10268 20532 10294 20535
rect 10268 20503 10294 20506
rect 10274 20093 10288 20503
rect 10406 20260 10432 20263
rect 10406 20231 10432 20234
rect 10268 20090 10294 20093
rect 10268 20061 10294 20064
rect 10274 20025 10288 20061
rect 10268 20022 10294 20025
rect 10268 19993 10294 19996
rect 10314 19920 10340 19923
rect 10314 19891 10340 19894
rect 10320 19719 10334 19891
rect 10314 19716 10340 19719
rect 10314 19687 10340 19690
rect 10360 19716 10386 19719
rect 10360 19687 10386 19690
rect 10366 18733 10380 19687
rect 10360 18730 10386 18733
rect 10360 18701 10386 18704
rect 10222 18424 10248 18427
rect 10222 18395 10248 18398
rect 10314 18390 10340 18393
rect 10314 18361 10340 18364
rect 10176 18288 10202 18291
rect 10176 18259 10202 18262
rect 10182 18087 10196 18259
rect 10320 18087 10334 18361
rect 10176 18084 10202 18087
rect 10176 18055 10202 18058
rect 10314 18084 10340 18087
rect 10314 18055 10340 18058
rect 10182 17237 10196 18055
rect 10412 18053 10426 20231
rect 10734 19753 10748 23325
rect 10866 23286 10892 23289
rect 10866 23257 10892 23260
rect 10872 23051 10886 23257
rect 10866 23048 10892 23051
rect 10866 23019 10892 23022
rect 10774 21552 10800 21555
rect 10774 21523 10800 21526
rect 10780 21351 10794 21523
rect 10774 21348 10800 21351
rect 10774 21319 10800 21322
rect 10820 21348 10846 21351
rect 10820 21319 10846 21322
rect 10728 19750 10754 19753
rect 10728 19721 10754 19724
rect 10774 18628 10800 18631
rect 10773 18612 10774 18616
rect 10800 18612 10801 18616
rect 10773 18579 10801 18584
rect 10780 18189 10794 18579
rect 10826 18412 10840 21319
rect 10872 21317 10886 23019
rect 11056 22983 11070 23555
rect 11378 23518 11392 24583
rect 11418 23524 11444 23527
rect 11378 23504 11418 23518
rect 11418 23495 11444 23498
rect 11424 22983 11438 23495
rect 11648 23286 11674 23289
rect 11648 23257 11674 23260
rect 11050 22980 11076 22983
rect 11050 22951 11076 22954
rect 11418 22980 11444 22983
rect 11444 22954 11484 22957
rect 11418 22951 11484 22954
rect 11424 22943 11484 22951
rect 11470 21895 11484 22943
rect 11556 22912 11582 22915
rect 11556 22883 11582 22886
rect 11562 22745 11576 22883
rect 11654 22813 11668 23257
rect 11648 22810 11674 22813
rect 11648 22781 11674 22784
rect 11556 22742 11582 22745
rect 11556 22713 11582 22716
rect 11555 22080 11583 22084
rect 11555 22047 11583 22052
rect 11372 21892 11398 21895
rect 11464 21892 11490 21895
rect 11398 21866 11438 21869
rect 11372 21863 11438 21866
rect 11464 21863 11490 21866
rect 11378 21855 11438 21863
rect 11424 21623 11438 21855
rect 11470 21657 11484 21863
rect 11562 21861 11576 22047
rect 11556 21858 11582 21861
rect 11556 21829 11582 21832
rect 11464 21654 11490 21657
rect 11464 21625 11490 21628
rect 11418 21620 11444 21623
rect 11418 21591 11444 21594
rect 11424 21351 11438 21591
rect 11050 21348 11076 21351
rect 11050 21319 11076 21322
rect 11418 21348 11444 21351
rect 11418 21319 11444 21322
rect 10866 21314 10892 21317
rect 10866 21285 10892 21288
rect 10958 21314 10984 21317
rect 10958 21285 10984 21288
rect 10964 21113 10978 21285
rect 11056 21283 11070 21319
rect 11470 21317 11484 21625
rect 11464 21314 11490 21317
rect 11464 21285 11490 21288
rect 11050 21280 11076 21283
rect 11050 21251 11076 21254
rect 10958 21110 10984 21113
rect 10958 21081 10984 21084
rect 10964 20807 10978 21081
rect 10958 20804 10984 20807
rect 10958 20775 10984 20778
rect 11056 20535 11070 21251
rect 11095 21128 11123 21132
rect 11095 21095 11123 21100
rect 11050 20532 11076 20535
rect 11050 20503 11076 20506
rect 11056 19821 11070 20503
rect 11050 19818 11076 19821
rect 11050 19789 11076 19792
rect 11050 18628 11076 18631
rect 11102 18622 11116 21095
rect 11234 20906 11260 20909
rect 11234 20877 11260 20880
rect 11280 20906 11306 20909
rect 11280 20877 11306 20880
rect 11141 20856 11169 20860
rect 11141 20823 11169 20828
rect 11148 20263 11162 20823
rect 11240 20781 11254 20877
rect 11286 20860 11300 20877
rect 11279 20856 11307 20860
rect 11279 20823 11307 20828
rect 11240 20767 11300 20781
rect 11286 20739 11300 20767
rect 11280 20736 11306 20739
rect 11280 20707 11306 20710
rect 11470 20569 11484 21285
rect 11562 21079 11576 21829
rect 11878 21688 11904 21691
rect 11878 21659 11904 21662
rect 11884 21472 11898 21659
rect 11877 21468 11905 21472
rect 11877 21435 11905 21440
rect 11648 21314 11674 21317
rect 11648 21285 11674 21288
rect 11556 21076 11582 21079
rect 11556 21047 11582 21050
rect 11654 20909 11668 21285
rect 11648 20906 11674 20909
rect 11648 20877 11674 20880
rect 11832 20804 11858 20807
rect 11832 20775 11858 20778
rect 11372 20566 11398 20569
rect 11372 20537 11398 20540
rect 11464 20566 11490 20569
rect 11464 20537 11490 20540
rect 11142 20260 11168 20263
rect 11142 20231 11168 20234
rect 11378 20229 11392 20537
rect 11418 20532 11444 20535
rect 11418 20503 11444 20506
rect 11424 20297 11438 20503
rect 11418 20294 11444 20297
rect 11418 20265 11444 20268
rect 11372 20226 11398 20229
rect 11372 20197 11398 20200
rect 11378 19719 11392 20197
rect 11786 20022 11812 20025
rect 11838 20016 11852 20775
rect 11884 20365 11898 21435
rect 11878 20362 11904 20365
rect 11878 20333 11904 20336
rect 11923 20040 11951 20044
rect 11812 20002 11852 20016
rect 11878 20022 11904 20025
rect 11786 19993 11812 19996
rect 11923 20007 11924 20012
rect 11878 19993 11904 19996
rect 11950 20007 11951 20012
rect 11924 19993 11950 19996
rect 11884 19821 11898 19993
rect 11878 19818 11904 19821
rect 11878 19789 11904 19792
rect 11372 19716 11398 19719
rect 11187 19700 11215 19704
rect 11372 19687 11398 19690
rect 11187 19667 11188 19672
rect 11214 19667 11215 19672
rect 11188 19653 11214 19656
rect 11194 19549 11208 19653
rect 11188 19546 11214 19549
rect 11188 19517 11214 19520
rect 11464 18934 11490 18937
rect 11464 18905 11490 18908
rect 11076 18608 11116 18622
rect 11050 18599 11076 18602
rect 11470 18597 11484 18905
rect 11832 18900 11858 18903
rect 11832 18871 11858 18874
rect 11838 18631 11852 18871
rect 11832 18628 11858 18631
rect 11832 18599 11858 18602
rect 10866 18594 10892 18597
rect 10866 18565 10892 18568
rect 11004 18594 11030 18597
rect 11004 18565 11030 18568
rect 11464 18594 11490 18597
rect 11464 18565 11490 18568
rect 11648 18594 11674 18597
rect 11648 18565 11674 18568
rect 10819 18408 10847 18412
rect 10819 18375 10847 18380
rect 10872 18189 10886 18565
rect 10912 18560 10938 18563
rect 10912 18531 10938 18534
rect 10774 18186 10800 18189
rect 10774 18157 10800 18160
rect 10866 18186 10892 18189
rect 10866 18157 10892 18160
rect 10406 18050 10432 18053
rect 10406 18021 10432 18024
rect 10918 17237 10932 18531
rect 11010 18461 11024 18565
rect 11654 18461 11668 18565
rect 11004 18458 11030 18461
rect 11004 18429 11030 18432
rect 11648 18458 11674 18461
rect 11648 18429 11674 18432
rect 11188 17472 11214 17475
rect 11188 17443 11214 17446
rect 10176 17234 10202 17237
rect 10176 17205 10202 17208
rect 10590 17234 10616 17237
rect 10590 17205 10616 17208
rect 10912 17234 10938 17237
rect 10912 17205 10938 17208
rect 10130 16962 10156 16965
rect 10130 16933 10156 16936
rect 10136 16769 10150 16933
rect 10136 16761 10196 16769
rect 9532 16758 9558 16761
rect 9532 16729 9558 16732
rect 9624 16758 9650 16761
rect 9624 16729 9650 16732
rect 9670 16758 9696 16761
rect 9670 16729 9696 16732
rect 10038 16758 10064 16761
rect 10136 16758 10202 16761
rect 10136 16755 10176 16758
rect 10038 16729 10064 16732
rect 10176 16729 10202 16732
rect 9676 16557 9690 16729
rect 9808 16656 9834 16659
rect 9808 16627 9834 16630
rect 9670 16554 9696 16557
rect 9670 16525 9696 16528
rect 9814 16455 9828 16627
rect 9854 16520 9880 16523
rect 9854 16491 9880 16494
rect 9808 16452 9834 16455
rect 9808 16423 9834 16426
rect 9348 15874 9374 15877
rect 9348 15845 9374 15848
rect 9256 15670 9282 15673
rect 9256 15641 9282 15644
rect 9210 15126 9236 15129
rect 9210 15097 9236 15100
rect 9164 15092 9190 15095
rect 9164 15063 9190 15066
rect 9118 15024 9144 15027
rect 9118 14995 9144 14998
rect 8934 14820 8960 14823
rect 8934 14791 8960 14794
rect 8980 14820 9006 14823
rect 8980 14791 9006 14794
rect 8888 14786 8914 14789
rect 8888 14757 8914 14760
rect 8940 14585 8954 14791
rect 8934 14582 8960 14585
rect 8934 14553 8960 14556
rect 8842 14378 8868 14381
rect 8842 14349 8868 14352
rect 8704 14276 8730 14279
rect 8704 14247 8730 14250
rect 8474 13766 8500 13769
rect 8474 13737 8500 13740
rect 8290 13528 8316 13531
rect 8290 13499 8316 13502
rect 8106 13426 8132 13429
rect 8106 13397 8132 13400
rect 8014 13392 8040 13395
rect 8014 13363 8040 13366
rect 8020 13191 8034 13363
rect 8112 13191 8126 13397
rect 8198 13290 8224 13293
rect 8198 13261 8224 13264
rect 8204 13244 8218 13261
rect 8296 13259 8310 13499
rect 8290 13256 8316 13259
rect 8197 13240 8225 13244
rect 8290 13227 8316 13230
rect 8197 13207 8225 13212
rect 8204 13191 8218 13207
rect 8480 13191 8494 13737
rect 8612 13732 8638 13735
rect 8888 13732 8914 13735
rect 8612 13703 8638 13706
rect 8749 13716 8777 13720
rect 7876 13188 7902 13191
rect 7876 13159 7902 13162
rect 7922 13188 7948 13191
rect 7922 13159 7948 13162
rect 8014 13188 8040 13191
rect 8014 13159 8040 13162
rect 8089 13188 8126 13191
rect 8115 13176 8126 13188
rect 8198 13188 8224 13191
rect 8115 13172 8133 13176
rect 8089 13159 8105 13162
rect 7232 12644 7258 12647
rect 7232 12615 7258 12618
rect 7416 12610 7442 12613
rect 7416 12581 7442 12584
rect 7140 12406 7166 12409
rect 7100 12386 7140 12400
rect 7100 11865 7114 12386
rect 7140 12377 7166 12380
rect 7422 12205 7436 12581
rect 7599 12424 7627 12428
rect 7882 12409 7896 13159
rect 7928 12428 7942 13159
rect 8198 13159 8224 13162
rect 8474 13188 8500 13191
rect 8474 13159 8500 13162
rect 8105 13139 8133 13144
rect 8152 13120 8178 13123
rect 8152 13091 8178 13094
rect 8158 13021 8172 13091
rect 8152 13018 8178 13021
rect 8152 12989 8178 12992
rect 8336 12746 8362 12749
rect 8336 12717 8362 12720
rect 8342 12613 8356 12717
rect 8152 12610 8178 12613
rect 8152 12581 8178 12584
rect 8336 12610 8362 12613
rect 8336 12581 8362 12584
rect 8158 12443 8172 12581
rect 8152 12440 8178 12443
rect 7921 12424 7949 12428
rect 7599 12391 7627 12396
rect 7876 12406 7902 12409
rect 7416 12202 7442 12205
rect 7416 12173 7442 12176
rect 7324 12100 7350 12103
rect 7324 12071 7350 12074
rect 7416 12100 7442 12103
rect 7416 12071 7442 12074
rect 7462 12100 7488 12103
rect 7462 12071 7488 12074
rect 7554 12100 7580 12103
rect 7606 12077 7620 12391
rect 8152 12411 8178 12414
rect 8480 12409 8494 13159
rect 8618 13157 8632 13703
rect 8940 13726 8954 14553
rect 9124 14551 9138 14995
rect 9118 14548 9144 14551
rect 9118 14519 9144 14522
rect 9170 14497 9184 15063
rect 9216 14925 9230 15097
rect 9210 14922 9236 14925
rect 9210 14893 9236 14896
rect 9262 14585 9276 15641
rect 9354 14619 9368 15845
rect 9348 14616 9374 14619
rect 9348 14587 9374 14590
rect 9256 14582 9282 14585
rect 9256 14553 9282 14556
rect 9032 14483 9184 14497
rect 9032 13807 9046 14483
rect 9624 14038 9650 14041
rect 9624 14009 9650 14012
rect 9762 14038 9788 14041
rect 9762 14009 9788 14012
rect 9630 13837 9644 14009
rect 9670 13936 9696 13939
rect 9670 13907 9696 13910
rect 8914 13712 8954 13726
rect 8986 13793 9046 13807
rect 9624 13834 9650 13837
rect 9624 13805 9650 13808
rect 8888 13703 8914 13706
rect 8749 13683 8750 13688
rect 8776 13683 8777 13688
rect 8750 13669 8776 13672
rect 8986 13380 9000 13793
rect 9676 13565 9690 13907
rect 9670 13562 9696 13565
rect 9670 13533 9696 13536
rect 9256 13494 9282 13497
rect 9256 13465 9282 13468
rect 8979 13376 9007 13380
rect 8979 13343 9007 13348
rect 8612 13154 8638 13157
rect 8612 13125 8638 13128
rect 8618 12443 8632 13125
rect 8612 12440 8638 12443
rect 8612 12411 8638 12414
rect 7921 12391 7949 12396
rect 8474 12406 8500 12409
rect 7876 12377 7902 12380
rect 8474 12377 8500 12380
rect 8480 12137 8494 12377
rect 8474 12134 8500 12137
rect 8474 12105 8500 12108
rect 7580 12074 7620 12077
rect 7554 12071 7620 12074
rect 7330 11952 7344 12071
rect 7323 11948 7351 11952
rect 7323 11915 7351 11920
rect 7330 11899 7344 11915
rect 7324 11896 7350 11899
rect 7324 11867 7350 11870
rect 7094 11862 7120 11865
rect 7094 11833 7120 11836
rect 7422 11661 7436 12071
rect 7416 11658 7442 11661
rect 7416 11629 7442 11632
rect 7468 11083 7482 12071
rect 7560 12063 7620 12071
rect 8480 11593 8494 12105
rect 8566 12066 8592 12069
rect 8618 12060 8632 12411
rect 8934 12304 8960 12307
rect 8934 12275 8960 12278
rect 8592 12046 8632 12060
rect 8566 12037 8592 12040
rect 8618 11865 8632 12046
rect 8796 12066 8822 12069
rect 8796 12037 8822 12040
rect 8612 11862 8638 11865
rect 8612 11833 8638 11836
rect 8474 11590 8500 11593
rect 8474 11561 8500 11564
rect 7600 11556 7626 11559
rect 7600 11527 7626 11530
rect 7554 11522 7580 11525
rect 7554 11493 7580 11496
rect 7560 11287 7574 11493
rect 7606 11389 7620 11527
rect 8618 11525 8632 11833
rect 8802 11816 8816 12037
rect 8940 11865 8954 12275
rect 8986 11865 9000 13343
rect 9118 12950 9144 12953
rect 9118 12921 9144 12924
rect 9026 12848 9052 12851
rect 9026 12819 9052 12822
rect 9032 12632 9046 12819
rect 9025 12628 9053 12632
rect 9124 12613 9138 12921
rect 9262 12749 9276 13465
rect 9768 13123 9782 14009
rect 9860 13531 9874 16491
rect 10596 16489 10610 17205
rect 10918 17033 10932 17205
rect 10912 17030 10938 17033
rect 10912 17001 10938 17004
rect 11194 16965 11208 17443
rect 11648 17200 11674 17203
rect 11648 17171 11674 17174
rect 10636 16962 10662 16965
rect 10636 16933 10662 16936
rect 11188 16962 11214 16965
rect 11188 16933 11214 16936
rect 10590 16486 10616 16489
rect 10590 16457 10616 16460
rect 10642 16387 10656 16933
rect 10268 16384 10294 16387
rect 10268 16355 10294 16358
rect 10636 16384 10662 16387
rect 10636 16355 10662 16358
rect 10274 16285 10288 16355
rect 10268 16282 10294 16285
rect 10268 16253 10294 16256
rect 10642 15843 10656 16355
rect 11194 16304 11208 16933
rect 11654 16795 11668 17171
rect 11976 17101 11990 26691
rect 12206 26349 12220 26759
rect 13126 26757 13140 27303
rect 13258 27264 13284 27267
rect 13258 27235 13284 27238
rect 13264 27063 13278 27235
rect 13310 27097 13324 27541
rect 13356 27165 13370 27609
rect 13402 27267 13416 27609
rect 13396 27264 13422 27267
rect 13396 27235 13422 27238
rect 13350 27162 13376 27165
rect 13350 27133 13376 27136
rect 13304 27094 13330 27097
rect 13304 27065 13330 27068
rect 13258 27060 13284 27063
rect 13258 27031 13284 27034
rect 13120 26754 13146 26757
rect 13120 26725 13146 26728
rect 12246 26720 12272 26723
rect 12246 26691 12272 26694
rect 12252 26587 12266 26691
rect 12246 26584 12272 26587
rect 12246 26555 12272 26558
rect 12476 26448 12502 26451
rect 12476 26419 12502 26422
rect 12200 26346 12226 26349
rect 12200 26317 12226 26320
rect 12482 26247 12496 26419
rect 13264 26247 13278 27031
rect 13586 27029 13600 27609
rect 13718 27060 13744 27063
rect 13718 27031 13744 27034
rect 13580 27026 13606 27029
rect 13580 26997 13606 27000
rect 13488 26550 13514 26553
rect 13488 26521 13514 26524
rect 13534 26550 13560 26553
rect 13534 26521 13560 26524
rect 12476 26244 12502 26247
rect 12476 26215 12502 26218
rect 13028 26244 13054 26247
rect 13028 26215 13054 26218
rect 13258 26244 13284 26247
rect 13258 26215 13284 26218
rect 12062 25088 12088 25091
rect 12062 25059 12088 25062
rect 12068 24377 12082 25059
rect 12430 24816 12456 24819
rect 12430 24787 12456 24790
rect 12338 24714 12364 24717
rect 12338 24685 12364 24688
rect 12154 24544 12180 24547
rect 12154 24515 12180 24518
rect 12108 24442 12134 24445
rect 12108 24413 12134 24416
rect 12016 24374 12042 24377
rect 12016 24345 12042 24348
rect 12062 24374 12088 24377
rect 12062 24345 12088 24348
rect 12022 24328 12036 24345
rect 12015 24324 12043 24328
rect 12015 24291 12043 24296
rect 12016 23456 12042 23459
rect 12016 23427 12042 23430
rect 12022 23323 12036 23427
rect 12114 23323 12128 24413
rect 12160 24377 12174 24515
rect 12344 24377 12358 24685
rect 12384 24646 12410 24649
rect 12384 24617 12410 24620
rect 12154 24374 12180 24377
rect 12154 24345 12180 24348
rect 12338 24374 12364 24377
rect 12338 24345 12364 24348
rect 12390 24309 12404 24617
rect 12436 24411 12450 24787
rect 12430 24408 12456 24411
rect 12430 24379 12456 24382
rect 12384 24306 12410 24309
rect 12384 24277 12410 24280
rect 12154 24272 12180 24275
rect 12154 24243 12180 24246
rect 12160 24071 12174 24243
rect 12154 24068 12180 24071
rect 12154 24039 12180 24042
rect 12292 24068 12318 24071
rect 12292 24039 12318 24042
rect 12016 23320 12042 23323
rect 12016 23291 12042 23294
rect 12108 23320 12134 23323
rect 12108 23291 12134 23294
rect 12114 23187 12128 23291
rect 12154 23286 12180 23289
rect 12154 23257 12180 23260
rect 12108 23184 12134 23187
rect 12108 23155 12134 23158
rect 12160 23085 12174 23257
rect 12298 23255 12312 24039
rect 12390 23629 12404 24277
rect 12384 23626 12410 23629
rect 12384 23597 12410 23600
rect 12292 23252 12318 23255
rect 12292 23223 12318 23226
rect 12154 23082 12180 23085
rect 12154 23053 12180 23056
rect 12430 21824 12456 21827
rect 12430 21795 12456 21798
rect 12338 21552 12364 21555
rect 12338 21523 12364 21526
rect 12344 21181 12358 21523
rect 12338 21178 12364 21181
rect 12338 21149 12364 21152
rect 12383 21128 12411 21132
rect 12436 21113 12450 21795
rect 12383 21095 12384 21100
rect 12410 21095 12411 21100
rect 12430 21110 12456 21113
rect 12384 21081 12410 21084
rect 12430 21081 12456 21084
rect 12384 20464 12410 20467
rect 12344 20444 12384 20458
rect 12016 20362 12042 20365
rect 12016 20333 12042 20336
rect 12022 20093 12036 20333
rect 12016 20090 12042 20093
rect 12016 20061 12042 20064
rect 12344 20025 12358 20444
rect 12384 20435 12410 20438
rect 12383 20244 12411 20248
rect 12383 20211 12411 20216
rect 12390 20025 12404 20211
rect 12430 20192 12456 20195
rect 12430 20163 12456 20166
rect 12436 20093 12450 20163
rect 12430 20090 12456 20093
rect 12430 20061 12456 20064
rect 12338 20022 12364 20025
rect 12338 19993 12364 19996
rect 12384 20022 12410 20025
rect 12482 20016 12496 26215
rect 13034 26009 13048 26215
rect 13264 26179 13278 26215
rect 13258 26176 13284 26179
rect 13258 26147 13284 26150
rect 13028 26006 13054 26009
rect 13028 25977 13054 25980
rect 13264 25941 13278 26147
rect 13120 25938 13146 25941
rect 13120 25909 13146 25912
rect 13258 25938 13284 25941
rect 13258 25909 13284 25912
rect 12982 25904 13008 25907
rect 12982 25875 13008 25878
rect 12988 25703 13002 25875
rect 12982 25700 13008 25703
rect 12982 25671 13008 25674
rect 12844 25258 12870 25261
rect 12844 25229 12870 25232
rect 12798 24918 12824 24921
rect 12798 24889 12824 24892
rect 12804 24547 12818 24889
rect 12798 24544 12824 24547
rect 12798 24515 12824 24518
rect 12660 24068 12686 24071
rect 12660 24039 12686 24042
rect 12666 21691 12680 24039
rect 12660 21688 12686 21691
rect 12660 21659 12686 21662
rect 12706 21654 12732 21657
rect 12706 21625 12732 21628
rect 12614 21552 12640 21555
rect 12614 21523 12640 21526
rect 12522 21280 12548 21283
rect 12522 21251 12548 21254
rect 12528 21113 12542 21251
rect 12522 21110 12548 21113
rect 12522 21081 12548 21084
rect 12620 21079 12634 21523
rect 12660 21178 12686 21181
rect 12660 21149 12686 21152
rect 12614 21076 12640 21079
rect 12614 21047 12640 21050
rect 12666 21045 12680 21149
rect 12660 21042 12686 21045
rect 12660 21013 12686 21016
rect 12568 20872 12594 20875
rect 12568 20843 12594 20846
rect 12384 19993 12410 19996
rect 12436 20002 12496 20016
rect 12062 19920 12088 19923
rect 12062 19891 12088 19894
rect 12068 19821 12082 19891
rect 12062 19818 12088 19821
rect 12062 19789 12088 19792
rect 12390 19379 12404 19993
rect 12384 19376 12410 19379
rect 12384 19347 12410 19350
rect 12108 19104 12134 19107
rect 12108 19075 12134 19078
rect 12114 18937 12128 19075
rect 12436 19013 12450 20002
rect 12522 19784 12548 19787
rect 12522 19755 12548 19758
rect 12528 19481 12542 19755
rect 12522 19478 12548 19481
rect 12522 19449 12548 19452
rect 12436 18999 12496 19013
rect 12108 18934 12134 18937
rect 12108 18905 12134 18908
rect 12430 18934 12456 18937
rect 12430 18905 12456 18908
rect 12436 17883 12450 18905
rect 12430 17880 12456 17883
rect 12430 17851 12456 17854
rect 11970 17098 11996 17101
rect 11970 17069 11996 17072
rect 12246 16996 12272 16999
rect 12245 16980 12246 16984
rect 12272 16980 12273 16984
rect 12245 16947 12273 16952
rect 12108 16928 12134 16931
rect 12108 16899 12134 16902
rect 11648 16792 11674 16795
rect 11648 16763 11674 16766
rect 11739 16776 11767 16780
rect 11694 16758 11720 16761
rect 12114 16761 12128 16899
rect 11739 16743 11740 16748
rect 11694 16729 11720 16732
rect 11766 16743 11767 16748
rect 12108 16758 12134 16761
rect 11740 16729 11766 16732
rect 12108 16729 12134 16732
rect 11700 16557 11714 16729
rect 11746 16659 11760 16729
rect 11740 16656 11766 16659
rect 11740 16627 11766 16630
rect 12154 16656 12180 16659
rect 12154 16627 12180 16630
rect 11694 16554 11720 16557
rect 11694 16525 11720 16528
rect 11187 16300 11215 16304
rect 11187 16267 11215 16272
rect 10774 15908 10800 15911
rect 10774 15879 10800 15882
rect 10636 15840 10662 15843
rect 10636 15811 10662 15814
rect 10452 15568 10478 15571
rect 10452 15539 10478 15542
rect 10268 15160 10294 15163
rect 10268 15131 10294 15134
rect 10176 15024 10202 15027
rect 10176 14995 10202 14998
rect 10182 14823 10196 14995
rect 10176 14820 10202 14823
rect 10176 14791 10202 14794
rect 10176 14752 10202 14755
rect 10176 14723 10202 14726
rect 10038 13732 10064 13735
rect 10038 13703 10064 13706
rect 9854 13528 9880 13531
rect 9854 13499 9880 13502
rect 10044 13463 10058 13703
rect 10038 13460 10064 13463
rect 10038 13431 10064 13434
rect 9946 13392 9972 13395
rect 9946 13363 9972 13366
rect 9762 13120 9788 13123
rect 9762 13091 9788 13094
rect 9256 12746 9282 12749
rect 9256 12717 9282 12720
rect 9025 12595 9053 12600
rect 9118 12610 9144 12613
rect 9032 12443 9046 12595
rect 9118 12581 9144 12584
rect 9026 12440 9052 12443
rect 9026 12411 9052 12414
rect 9669 12152 9697 12156
rect 9669 12119 9697 12124
rect 9118 12100 9144 12103
rect 9118 12071 9144 12074
rect 9124 11884 9138 12071
rect 9532 12032 9558 12035
rect 9532 12003 9558 12006
rect 9117 11880 9145 11884
rect 8934 11862 8960 11865
rect 8934 11833 8960 11836
rect 8980 11862 9006 11865
rect 9538 11865 9552 12003
rect 9676 11865 9690 12119
rect 9716 11896 9742 11899
rect 9716 11867 9742 11870
rect 9117 11847 9118 11852
rect 8980 11833 9006 11836
rect 9144 11847 9145 11852
rect 9532 11862 9558 11865
rect 9118 11833 9144 11836
rect 9532 11833 9558 11836
rect 9578 11862 9604 11865
rect 9578 11833 9604 11836
rect 9670 11862 9696 11865
rect 9670 11833 9696 11836
rect 8795 11812 8823 11816
rect 8795 11779 8823 11784
rect 9584 11748 9598 11833
rect 9577 11744 9605 11748
rect 9577 11711 9605 11716
rect 9584 11661 9598 11711
rect 9578 11658 9604 11661
rect 9578 11629 9604 11632
rect 8704 11556 8730 11559
rect 8704 11527 8730 11530
rect 8612 11522 8638 11525
rect 8612 11493 8638 11496
rect 8710 11476 8724 11527
rect 8703 11472 8731 11476
rect 8703 11439 8731 11444
rect 9676 11389 9690 11833
rect 9722 11661 9736 11867
rect 9900 11828 9926 11831
rect 9900 11799 9926 11802
rect 9716 11658 9742 11661
rect 9716 11629 9742 11632
rect 9906 11559 9920 11799
rect 9900 11556 9926 11559
rect 9900 11527 9926 11530
rect 9952 11525 9966 13363
rect 10044 13225 10058 13431
rect 10083 13308 10111 13312
rect 10083 13275 10084 13280
rect 10110 13275 10111 13280
rect 10084 13261 10110 13264
rect 10038 13222 10064 13225
rect 10038 13193 10064 13196
rect 10044 12919 10058 13193
rect 10090 12987 10104 13261
rect 10084 12984 10110 12987
rect 10084 12955 10110 12958
rect 10038 12916 10064 12919
rect 10038 12887 10064 12890
rect 10044 12681 10058 12887
rect 10038 12678 10064 12681
rect 10038 12649 10064 12652
rect 10044 12409 10058 12649
rect 10038 12406 10064 12409
rect 10038 12377 10064 12380
rect 10044 12137 10058 12377
rect 10038 12134 10064 12137
rect 10038 12105 10064 12108
rect 9991 11948 10019 11952
rect 9991 11915 10019 11920
rect 9998 11899 10012 11915
rect 9992 11896 10018 11899
rect 9992 11867 10018 11870
rect 10182 11593 10196 14723
rect 10274 14619 10288 15131
rect 10458 14891 10472 15539
rect 10780 15401 10794 15879
rect 10820 15874 10846 15877
rect 10820 15845 10846 15848
rect 10774 15398 10800 15401
rect 10774 15369 10800 15372
rect 10544 15194 10570 15197
rect 10544 15165 10570 15168
rect 10452 14888 10478 14891
rect 10452 14859 10478 14862
rect 10550 14789 10564 15165
rect 10780 14857 10794 15369
rect 10826 15358 10840 15845
rect 11832 15840 11858 15843
rect 11832 15811 11858 15814
rect 11096 15704 11122 15707
rect 11096 15675 11122 15678
rect 10912 15364 10938 15367
rect 10826 15344 10912 15358
rect 10912 15335 10938 15338
rect 10918 15129 10932 15335
rect 11102 15333 11116 15675
rect 11142 15364 11168 15367
rect 11142 15335 11168 15338
rect 11096 15330 11122 15333
rect 11096 15301 11122 15304
rect 10912 15126 10938 15129
rect 10912 15097 10938 15100
rect 10774 14854 10800 14857
rect 10774 14825 10800 14828
rect 10544 14786 10570 14789
rect 10544 14757 10570 14760
rect 10360 14752 10386 14755
rect 10360 14723 10386 14726
rect 10268 14616 10294 14619
rect 10268 14587 10294 14590
rect 10366 14483 10380 14723
rect 10360 14480 10386 14483
rect 10360 14451 10386 14454
rect 10780 14279 10794 14825
rect 11148 14279 11162 15335
rect 11838 15129 11852 15811
rect 11970 15296 11996 15299
rect 11970 15267 11996 15270
rect 11976 15197 11990 15267
rect 11970 15194 11996 15197
rect 11970 15165 11996 15168
rect 12107 15144 12135 15148
rect 11832 15126 11858 15129
rect 11832 15097 11858 15100
rect 12062 15126 12088 15129
rect 12107 15111 12135 15116
rect 12062 15097 12088 15100
rect 12016 15024 12042 15027
rect 12016 14995 12042 14998
rect 11418 14854 11444 14857
rect 11418 14825 11444 14828
rect 11424 14585 11438 14825
rect 11694 14820 11720 14823
rect 11694 14791 11720 14794
rect 11740 14820 11766 14823
rect 11740 14791 11766 14794
rect 11700 14653 11714 14791
rect 11694 14650 11720 14653
rect 11694 14621 11720 14624
rect 11746 14619 11760 14791
rect 11740 14616 11766 14619
rect 11740 14587 11766 14590
rect 11418 14582 11444 14585
rect 11418 14553 11444 14556
rect 10774 14276 10800 14279
rect 10774 14247 10800 14250
rect 11004 14276 11030 14279
rect 11004 14247 11030 14250
rect 11142 14276 11168 14279
rect 11142 14247 11168 14250
rect 10780 13837 10794 14247
rect 10774 13834 10800 13837
rect 10774 13805 10800 13808
rect 11010 13735 11024 14247
rect 11096 14242 11122 14245
rect 11096 14213 11122 14216
rect 11102 14109 11116 14213
rect 11096 14106 11122 14109
rect 11096 14077 11122 14080
rect 11102 13777 11116 14077
rect 11056 13763 11116 13777
rect 10728 13732 10754 13735
rect 11004 13732 11030 13735
rect 10728 13703 10754 13706
rect 10911 13716 10939 13720
rect 10267 13580 10295 13584
rect 10267 13547 10295 13552
rect 10274 13531 10288 13547
rect 10268 13528 10294 13531
rect 10268 13499 10294 13502
rect 10274 12851 10288 13499
rect 10734 13497 10748 13703
rect 11004 13703 11030 13706
rect 10911 13683 10912 13688
rect 10938 13683 10939 13688
rect 10912 13669 10938 13672
rect 10314 13494 10340 13497
rect 10314 13465 10340 13468
rect 10728 13494 10754 13497
rect 10728 13465 10754 13468
rect 10320 12953 10334 13465
rect 11010 13157 11024 13703
rect 11056 13191 11070 13763
rect 11648 13528 11674 13531
rect 11648 13499 11674 13502
rect 11050 13188 11076 13191
rect 11050 13159 11076 13162
rect 11654 13157 11668 13499
rect 11878 13392 11904 13395
rect 11878 13363 11904 13366
rect 11739 13308 11767 13312
rect 11739 13275 11767 13280
rect 11746 13176 11760 13275
rect 11739 13172 11767 13176
rect 11004 13154 11030 13157
rect 11004 13125 11030 13128
rect 11280 13154 11306 13157
rect 11280 13125 11306 13128
rect 11648 13154 11674 13157
rect 11739 13139 11767 13144
rect 11648 13125 11674 13128
rect 10314 12950 10340 12953
rect 10314 12921 10340 12924
rect 10268 12848 10294 12851
rect 10268 12819 10294 12822
rect 10320 12647 10334 12921
rect 11286 12749 11300 13125
rect 11746 12953 11760 13139
rect 11884 12953 11898 13363
rect 11740 12950 11766 12953
rect 11740 12921 11766 12924
rect 11878 12950 11904 12953
rect 11878 12921 11904 12924
rect 11280 12746 11306 12749
rect 11280 12717 11306 12720
rect 10314 12644 10340 12647
rect 10314 12615 10340 12618
rect 10452 12644 10478 12647
rect 10452 12615 10478 12618
rect 10405 12492 10433 12496
rect 10405 12459 10406 12464
rect 10432 12459 10433 12464
rect 10406 12445 10432 12448
rect 10222 12100 10248 12103
rect 10222 12071 10248 12074
rect 10228 11865 10242 12071
rect 10412 12069 10426 12445
rect 10458 12103 10472 12615
rect 11694 12576 11720 12579
rect 11694 12547 11720 12550
rect 11700 12477 11714 12547
rect 11694 12474 11720 12477
rect 11694 12445 11720 12448
rect 12022 12443 12036 14995
rect 12068 14925 12082 15097
rect 12114 15095 12128 15111
rect 12108 15092 12134 15095
rect 12108 15063 12134 15066
rect 12062 14922 12088 14925
rect 12062 14893 12088 14896
rect 12160 14279 12174 16627
rect 12252 16523 12266 16947
rect 12292 16792 12318 16795
rect 12292 16763 12318 16766
rect 12246 16520 12272 16523
rect 12246 16491 12272 16494
rect 12298 14891 12312 16763
rect 12482 16557 12496 18999
rect 12574 18937 12588 20843
rect 12614 20736 12640 20739
rect 12614 20707 12640 20710
rect 12620 20059 12634 20707
rect 12614 20056 12640 20059
rect 12614 20027 12640 20030
rect 12614 19988 12640 19991
rect 12613 19972 12614 19976
rect 12640 19972 12641 19976
rect 12613 19939 12641 19944
rect 12620 19787 12634 19939
rect 12614 19784 12640 19787
rect 12614 19755 12640 19758
rect 12614 19546 12640 19549
rect 12614 19517 12640 19520
rect 12568 18934 12594 18937
rect 12568 18905 12594 18908
rect 12620 18877 12634 19517
rect 12574 18863 12634 18877
rect 12476 16554 12502 16557
rect 12476 16525 12502 16528
rect 12482 15877 12496 16525
rect 12482 15863 12542 15877
rect 12528 15673 12542 15863
rect 12522 15670 12548 15673
rect 12522 15641 12548 15644
rect 12384 15636 12410 15639
rect 12384 15607 12410 15610
rect 12390 15095 12404 15607
rect 12384 15092 12410 15095
rect 12384 15063 12410 15066
rect 12292 14888 12318 14891
rect 12292 14859 12318 14862
rect 12292 14820 12318 14823
rect 12318 14800 12358 14814
rect 12292 14791 12318 14794
rect 12154 14276 12180 14279
rect 12154 14247 12180 14250
rect 12200 14276 12226 14279
rect 12200 14247 12226 14250
rect 12206 13837 12220 14247
rect 12292 14242 12318 14245
rect 12292 14213 12318 14216
rect 12246 14208 12272 14211
rect 12246 14179 12272 14182
rect 12200 13834 12226 13837
rect 12200 13805 12226 13808
rect 12061 13240 12089 13244
rect 12061 13207 12089 13212
rect 12068 12953 12082 13207
rect 12252 12953 12266 14179
rect 12298 14075 12312 14213
rect 12344 14211 12358 14800
rect 12390 14585 12404 15063
rect 12528 14585 12542 15641
rect 12574 14925 12588 18863
rect 12666 18616 12680 21013
rect 12712 19957 12726 21625
rect 12752 21110 12778 21113
rect 12752 21081 12778 21084
rect 12758 20365 12772 21081
rect 12804 20875 12818 24515
rect 12850 23255 12864 25229
rect 12988 24615 13002 25671
rect 13126 24921 13140 25909
rect 13494 25703 13508 26521
rect 13540 26281 13554 26521
rect 13586 26519 13600 26997
rect 13626 26822 13652 26825
rect 13626 26793 13652 26796
rect 13632 26757 13646 26793
rect 13626 26754 13652 26757
rect 13626 26725 13652 26728
rect 13580 26516 13606 26519
rect 13580 26487 13606 26490
rect 13534 26278 13560 26281
rect 13534 26249 13560 26252
rect 13488 25700 13514 25703
rect 13488 25671 13514 25674
rect 13540 25669 13554 26249
rect 13586 25975 13600 26487
rect 13632 26281 13646 26725
rect 13672 26448 13698 26451
rect 13672 26419 13698 26422
rect 13626 26278 13652 26281
rect 13626 26249 13652 26252
rect 13678 26247 13692 26419
rect 13672 26244 13698 26247
rect 13672 26215 13698 26218
rect 13724 25975 13738 27031
rect 13764 26550 13790 26553
rect 13764 26521 13790 26524
rect 13770 26077 13784 26521
rect 13764 26074 13790 26077
rect 13764 26045 13790 26048
rect 13580 25972 13606 25975
rect 13580 25943 13606 25946
rect 13718 25972 13744 25975
rect 13718 25943 13744 25946
rect 13534 25666 13560 25669
rect 13534 25637 13560 25640
rect 13120 24918 13146 24921
rect 13120 24889 13146 24892
rect 13258 24918 13284 24921
rect 13258 24889 13284 24892
rect 12982 24612 13008 24615
rect 12982 24583 13008 24586
rect 12988 23527 13002 24583
rect 13212 24170 13238 24173
rect 13212 24141 13238 24144
rect 13120 23864 13146 23867
rect 13120 23835 13146 23838
rect 12982 23524 13008 23527
rect 12982 23495 13008 23498
rect 12890 23456 12916 23459
rect 12890 23427 12916 23430
rect 12844 23252 12870 23255
rect 12844 23223 12870 23226
rect 12798 20872 12824 20875
rect 12798 20843 12824 20846
rect 12798 20532 12824 20535
rect 12798 20503 12824 20506
rect 12752 20362 12778 20365
rect 12752 20333 12778 20336
rect 12752 20294 12778 20297
rect 12752 20265 12778 20268
rect 12758 19991 12772 20265
rect 12804 20263 12818 20503
rect 12798 20260 12824 20263
rect 12798 20231 12824 20234
rect 12752 19988 12778 19991
rect 12752 19959 12778 19962
rect 12706 19954 12732 19957
rect 12706 19925 12732 19928
rect 12758 19719 12772 19959
rect 12752 19716 12778 19719
rect 12752 19687 12778 19690
rect 12659 18612 12687 18616
rect 12659 18579 12687 18584
rect 12758 18359 12772 19687
rect 12804 18427 12818 20231
rect 12850 18461 12864 23223
rect 12896 21812 12910 23427
rect 12988 22745 13002 23495
rect 13126 23289 13140 23835
rect 13120 23286 13146 23289
rect 13120 23257 13146 23260
rect 13126 22983 13140 23257
rect 13120 22980 13146 22983
rect 13120 22951 13146 22954
rect 12982 22742 13008 22745
rect 12982 22713 13008 22716
rect 13028 22674 13054 22677
rect 13028 22645 13054 22648
rect 12889 21808 12917 21812
rect 12889 21775 12917 21780
rect 12844 18458 12870 18461
rect 12844 18429 12870 18432
rect 12798 18424 12824 18427
rect 12798 18395 12824 18398
rect 12752 18356 12778 18359
rect 12752 18327 12778 18330
rect 12758 18087 12772 18327
rect 12752 18084 12778 18087
rect 12752 18055 12778 18058
rect 12758 17849 12772 18055
rect 12752 17846 12778 17849
rect 12752 17817 12778 17820
rect 12614 17336 12640 17339
rect 12758 17313 12772 17817
rect 12614 17307 12640 17310
rect 12568 14922 12594 14925
rect 12568 14893 12594 14896
rect 12384 14582 12410 14585
rect 12384 14553 12410 14556
rect 12522 14582 12548 14585
rect 12522 14553 12548 14556
rect 12390 14536 12404 14553
rect 12383 14532 12411 14536
rect 12383 14499 12411 14504
rect 12384 14276 12410 14279
rect 12384 14247 12410 14250
rect 12338 14208 12364 14211
rect 12338 14179 12364 14182
rect 12292 14072 12318 14075
rect 12292 14043 12318 14046
rect 12390 13973 12404 14247
rect 12384 13970 12410 13973
rect 12384 13941 12410 13944
rect 12528 13497 12542 14553
rect 12430 13494 12456 13497
rect 12430 13465 12456 13468
rect 12522 13494 12548 13497
rect 12522 13465 12548 13468
rect 12436 13293 12450 13465
rect 12476 13392 12502 13395
rect 12476 13363 12502 13366
rect 12430 13290 12456 13293
rect 12430 13261 12456 13264
rect 12384 13018 12410 13021
rect 12384 12989 12410 12992
rect 12062 12950 12088 12953
rect 12062 12921 12088 12924
rect 12246 12950 12272 12953
rect 12246 12921 12272 12924
rect 12062 12882 12088 12885
rect 12062 12853 12088 12856
rect 12068 12749 12082 12853
rect 12062 12746 12088 12749
rect 12062 12717 12088 12720
rect 12390 12477 12404 12989
rect 12482 12953 12496 13363
rect 12476 12950 12502 12953
rect 12476 12921 12502 12924
rect 12430 12848 12456 12851
rect 12430 12819 12456 12822
rect 12384 12474 12410 12477
rect 12384 12445 12410 12448
rect 12016 12440 12042 12443
rect 11647 12424 11675 12428
rect 11556 12406 11582 12409
rect 12016 12411 12042 12414
rect 11647 12391 11648 12396
rect 11556 12377 11582 12380
rect 11674 12391 11675 12396
rect 11694 12406 11720 12409
rect 11648 12377 11674 12380
rect 11694 12377 11720 12380
rect 11740 12406 11766 12409
rect 11740 12377 11766 12380
rect 10866 12372 10892 12375
rect 10866 12343 10892 12346
rect 10452 12100 10478 12103
rect 10452 12071 10478 12074
rect 10406 12066 10432 12069
rect 10406 12037 10432 12040
rect 10222 11862 10248 11865
rect 10222 11833 10248 11836
rect 10458 11593 10472 12071
rect 10872 11831 10886 12343
rect 11562 12205 11576 12377
rect 11556 12202 11582 12205
rect 11556 12173 11582 12176
rect 11700 11933 11714 12377
rect 11694 11930 11720 11933
rect 11694 11901 11720 11904
rect 11746 11884 11760 12377
rect 11970 12304 11996 12307
rect 11970 12275 11996 12278
rect 11976 12137 11990 12275
rect 12015 12152 12043 12156
rect 11970 12134 11996 12137
rect 12015 12119 12043 12124
rect 11970 12105 11996 12108
rect 12022 12103 12036 12119
rect 12016 12100 12042 12103
rect 12016 12071 12042 12074
rect 11832 12066 11858 12069
rect 11832 12037 11858 12040
rect 11924 12066 11950 12069
rect 11924 12037 11950 12040
rect 11970 12066 11996 12069
rect 11970 12037 11996 12040
rect 11739 11880 11767 11884
rect 11739 11847 11767 11852
rect 10866 11828 10892 11831
rect 10866 11799 10892 11802
rect 11049 11812 11077 11816
rect 10872 11763 10886 11799
rect 11049 11779 11077 11784
rect 11647 11812 11675 11816
rect 11647 11779 11675 11784
rect 10866 11760 10892 11763
rect 10866 11731 10892 11734
rect 10176 11590 10202 11593
rect 10176 11561 10202 11564
rect 10452 11590 10478 11593
rect 10452 11561 10478 11564
rect 10872 11559 10886 11731
rect 10866 11556 10892 11559
rect 10866 11527 10892 11530
rect 9946 11522 9972 11525
rect 9946 11493 9972 11496
rect 10314 11488 10340 11491
rect 10314 11459 10340 11462
rect 7600 11386 7626 11389
rect 7600 11357 7626 11360
rect 9670 11386 9696 11389
rect 9670 11357 9696 11360
rect 7554 11284 7580 11287
rect 7554 11255 7580 11258
rect 7462 11080 7488 11083
rect 7462 11051 7488 11054
rect 5760 11012 5786 11015
rect 5760 10983 5786 10986
rect 6910 11012 6936 11015
rect 6910 10983 6936 10986
rect 10038 11012 10064 11015
rect 10038 10983 10064 10986
rect 10044 10777 10058 10983
rect 10320 10777 10334 11459
rect 10872 11015 10886 11527
rect 10866 11012 10892 11015
rect 10866 10983 10892 10986
rect 11056 10981 11070 11779
rect 11654 11661 11668 11779
rect 11648 11658 11674 11661
rect 11648 11629 11674 11632
rect 11096 11556 11122 11559
rect 11096 11527 11122 11530
rect 11102 11015 11116 11527
rect 11838 11049 11852 12037
rect 11930 11748 11944 12037
rect 11923 11744 11951 11748
rect 11923 11711 11951 11716
rect 11976 11661 11990 12037
rect 12384 11828 12410 11831
rect 12384 11799 12410 11802
rect 11970 11658 11996 11661
rect 11970 11629 11996 11632
rect 11832 11046 11858 11049
rect 11832 11017 11858 11020
rect 11096 11012 11122 11015
rect 11096 10983 11122 10986
rect 11050 10978 11076 10981
rect 11050 10949 11076 10952
rect 10038 10774 10064 10777
rect 10038 10745 10064 10748
rect 10314 10774 10340 10777
rect 10314 10745 10340 10748
rect 12390 10743 12404 11799
rect 12436 10811 12450 12819
rect 12620 12579 12634 17307
rect 12666 17305 12772 17313
rect 12660 17302 12772 17305
rect 12686 17299 12772 17302
rect 12660 17273 12686 17276
rect 12758 17033 12772 17299
rect 12752 17030 12778 17033
rect 12752 17001 12778 17004
rect 12660 16792 12686 16795
rect 12660 16763 12686 16766
rect 12666 14619 12680 16763
rect 12758 16761 12772 17001
rect 12752 16758 12778 16761
rect 12752 16729 12778 16732
rect 12758 16489 12772 16729
rect 12804 16659 12818 18395
rect 12850 17339 12864 18429
rect 12844 17336 12870 17339
rect 12844 17307 12870 17310
rect 12896 17052 12910 21775
rect 12982 21450 13008 21453
rect 12982 21421 13008 21424
rect 12988 21147 13002 21421
rect 12982 21144 13008 21147
rect 12935 21128 12963 21132
rect 12982 21115 13008 21118
rect 12935 21095 12936 21100
rect 12962 21095 12963 21100
rect 12936 21081 12962 21084
rect 12936 20838 12962 20841
rect 12936 20809 12962 20812
rect 12942 20297 12956 20809
rect 13034 20773 13048 22645
rect 13074 21654 13100 21657
rect 13074 21625 13100 21628
rect 13080 21351 13094 21625
rect 13074 21348 13100 21351
rect 13074 21319 13100 21322
rect 13074 21178 13100 21181
rect 13074 21149 13100 21152
rect 13080 20909 13094 21149
rect 13074 20906 13100 20909
rect 13074 20877 13100 20880
rect 13028 20770 13054 20773
rect 13028 20741 13054 20744
rect 13034 20535 13048 20741
rect 13074 20736 13100 20739
rect 13074 20707 13100 20710
rect 13028 20532 13054 20535
rect 13028 20503 13054 20506
rect 13028 20464 13054 20467
rect 13028 20435 13054 20438
rect 12936 20294 12962 20297
rect 12936 20265 12962 20268
rect 13034 20059 13048 20435
rect 13080 20263 13094 20707
rect 13074 20260 13100 20263
rect 13074 20231 13100 20234
rect 13028 20056 13054 20059
rect 13028 20027 13054 20030
rect 13080 19761 13094 20231
rect 13166 20226 13192 20229
rect 13166 20197 13192 20200
rect 13120 20022 13146 20025
rect 13120 19993 13146 19996
rect 13126 19976 13140 19993
rect 13119 19972 13147 19976
rect 13119 19939 13147 19944
rect 12988 19747 13094 19761
rect 12988 19651 13002 19747
rect 13028 19716 13054 19719
rect 13028 19687 13054 19690
rect 12982 19648 13008 19651
rect 12982 19619 13008 19622
rect 12988 19107 13002 19619
rect 12982 19104 13008 19107
rect 12982 19075 13008 19078
rect 12988 18699 13002 19075
rect 12982 18696 13008 18699
rect 12982 18667 13008 18670
rect 12936 18050 12962 18053
rect 12936 18021 12962 18024
rect 12942 17849 12956 18021
rect 12936 17846 12962 17849
rect 12936 17817 12962 17820
rect 12942 17305 12956 17817
rect 12936 17302 12962 17305
rect 12936 17273 12962 17276
rect 12889 17048 12917 17052
rect 12889 17015 12917 17020
rect 12844 16758 12870 16761
rect 12844 16729 12870 16732
rect 12798 16656 12824 16659
rect 12798 16627 12824 16630
rect 12752 16486 12778 16489
rect 12752 16457 12778 16460
rect 12758 16217 12772 16457
rect 12850 16217 12864 16729
rect 12896 16293 12910 17015
rect 12942 16965 12956 17273
rect 12936 16962 12962 16965
rect 12936 16933 12962 16936
rect 12942 16761 12956 16933
rect 13034 16795 13048 19687
rect 13172 19549 13186 20197
rect 13166 19546 13192 19549
rect 13166 19517 13192 19520
rect 13074 18832 13100 18835
rect 13074 18803 13100 18806
rect 13080 18631 13094 18803
rect 13074 18628 13100 18631
rect 13120 18628 13146 18631
rect 13074 18599 13100 18602
rect 13119 18612 13120 18616
rect 13146 18612 13147 18616
rect 13119 18579 13147 18584
rect 13074 18390 13100 18393
rect 13074 18361 13100 18364
rect 13080 18053 13094 18361
rect 13074 18050 13100 18053
rect 13074 18021 13100 18024
rect 13074 17880 13100 17883
rect 13074 17851 13100 17854
rect 13028 16792 13054 16795
rect 13028 16763 13054 16766
rect 12936 16758 12962 16761
rect 12936 16729 12962 16732
rect 13080 16701 13094 17851
rect 13166 16962 13192 16965
rect 13218 16956 13232 24141
rect 13264 23833 13278 24889
rect 13540 23867 13554 25637
rect 13810 24850 13836 24853
rect 13810 24821 13836 24824
rect 13816 24615 13830 24821
rect 13810 24612 13836 24615
rect 13810 24583 13836 24586
rect 13672 24544 13698 24547
rect 13672 24515 13698 24518
rect 13678 24173 13692 24515
rect 13816 24343 13830 24583
rect 13810 24340 13836 24343
rect 13810 24311 13836 24314
rect 13855 24324 13883 24328
rect 13855 24291 13883 24296
rect 13672 24170 13698 24173
rect 13672 24141 13698 24144
rect 13534 23864 13560 23867
rect 13534 23835 13560 23838
rect 13258 23830 13284 23833
rect 13258 23801 13284 23804
rect 13264 23527 13278 23801
rect 13304 23796 13330 23799
rect 13304 23767 13330 23770
rect 13258 23524 13284 23527
rect 13258 23495 13284 23498
rect 13258 23286 13284 23289
rect 13258 23257 13284 23260
rect 13264 22745 13278 23257
rect 13258 22742 13284 22745
rect 13258 22713 13284 22716
rect 13310 20807 13324 23767
rect 13396 22980 13422 22983
rect 13396 22951 13422 22954
rect 13402 22439 13416 22951
rect 13718 22742 13744 22745
rect 13718 22713 13744 22716
rect 13626 22674 13652 22677
rect 13626 22645 13652 22648
rect 13396 22436 13422 22439
rect 13396 22407 13422 22410
rect 13442 22368 13468 22371
rect 13442 22339 13468 22342
rect 13304 20804 13330 20807
rect 13304 20775 13330 20778
rect 13310 19719 13324 20775
rect 13448 20467 13462 22339
rect 13442 20464 13468 20467
rect 13442 20435 13468 20438
rect 13632 20263 13646 22645
rect 13724 22439 13738 22713
rect 13718 22436 13744 22439
rect 13718 22407 13744 22410
rect 13862 22371 13876 24291
rect 13902 24000 13928 24003
rect 13902 23971 13928 23974
rect 13908 23512 13922 23971
rect 13901 23508 13929 23512
rect 13901 23475 13929 23480
rect 13856 22368 13882 22371
rect 13856 22339 13882 22342
rect 13764 21314 13790 21317
rect 13764 21285 13790 21288
rect 13770 20773 13784 21285
rect 13764 20770 13790 20773
rect 13764 20741 13790 20744
rect 13626 20260 13652 20263
rect 13626 20231 13652 20234
rect 13304 19716 13330 19719
rect 13304 19687 13330 19690
rect 13672 18662 13698 18665
rect 13672 18633 13698 18636
rect 13678 18393 13692 18633
rect 13856 18628 13882 18631
rect 13856 18599 13882 18602
rect 13672 18390 13698 18393
rect 13672 18361 13698 18364
rect 13862 18189 13876 18599
rect 13856 18186 13882 18189
rect 13856 18157 13882 18160
rect 13625 18136 13653 18140
rect 13625 18103 13653 18108
rect 13632 18053 13646 18103
rect 13626 18050 13652 18053
rect 13626 18021 13652 18024
rect 13192 16942 13232 16956
rect 13166 16933 13192 16936
rect 13172 16848 13186 16933
rect 13165 16844 13193 16848
rect 13165 16811 13193 16816
rect 12988 16687 13094 16701
rect 12896 16279 12956 16293
rect 12942 16251 12956 16279
rect 12936 16248 12962 16251
rect 12936 16219 12962 16222
rect 12752 16214 12778 16217
rect 12752 16185 12778 16188
rect 12844 16214 12870 16217
rect 12844 16185 12870 16188
rect 12850 15163 12864 16185
rect 12844 15160 12870 15163
rect 12844 15131 12870 15134
rect 12660 14616 12686 14619
rect 12660 14587 12686 14590
rect 12936 13698 12962 13701
rect 12936 13669 12962 13672
rect 12942 13497 12956 13669
rect 12936 13494 12962 13497
rect 12936 13465 12962 13468
rect 12752 13460 12778 13463
rect 12752 13431 12778 13434
rect 12798 13460 12824 13463
rect 12798 13431 12824 13434
rect 12758 13293 12772 13431
rect 12752 13290 12778 13293
rect 12752 13261 12778 13264
rect 12804 13191 12818 13431
rect 12798 13188 12824 13191
rect 12798 13159 12824 13162
rect 12804 12919 12818 13159
rect 12942 13157 12956 13465
rect 12936 13154 12962 13157
rect 12936 13125 12962 13128
rect 12942 12953 12956 13125
rect 12988 13029 13002 16687
rect 13028 16656 13054 16659
rect 13028 16627 13054 16630
rect 13034 15673 13048 16627
rect 13172 16455 13186 16811
rect 13166 16452 13192 16455
rect 13166 16423 13192 16426
rect 13632 15877 13646 18021
rect 13908 17475 13922 23475
rect 13954 18087 13968 29173
rect 14086 28964 14112 28967
rect 14086 28935 14112 28938
rect 14092 28695 14106 28935
rect 14230 28748 14244 32968
rect 14322 32953 14336 32968
rect 14368 32953 14382 33000
rect 14322 32939 14382 32953
rect 15880 29814 15906 29817
rect 15880 29785 15906 29788
rect 15420 29576 15446 29579
rect 15420 29547 15446 29550
rect 15190 29304 15216 29307
rect 15190 29275 15216 29278
rect 14316 29270 14342 29273
rect 14316 29241 14342 29244
rect 14322 28899 14336 29241
rect 15006 29236 15032 29239
rect 15006 29207 15032 29210
rect 15012 29171 15026 29207
rect 15006 29168 15032 29171
rect 15006 29139 15032 29142
rect 15012 29035 15026 29139
rect 15196 29069 15210 29275
rect 15190 29066 15216 29069
rect 15190 29037 15216 29040
rect 15006 29032 15032 29035
rect 15006 29003 15032 29006
rect 15426 29001 15440 29547
rect 15696 29474 15722 29477
rect 15696 29445 15722 29448
rect 15702 29341 15716 29445
rect 15788 29440 15814 29443
rect 15788 29411 15814 29414
rect 15794 29341 15808 29411
rect 15696 29338 15722 29341
rect 15696 29309 15722 29312
rect 15788 29338 15814 29341
rect 15788 29309 15814 29312
rect 15794 29273 15808 29309
rect 15788 29270 15814 29273
rect 15788 29241 15814 29244
rect 15696 29032 15722 29035
rect 15696 29003 15722 29006
rect 15420 28998 15446 29001
rect 15420 28969 15446 28972
rect 14316 28896 14342 28899
rect 14316 28867 14342 28870
rect 14592 28896 14618 28899
rect 14592 28867 14618 28870
rect 14223 28744 14251 28748
rect 14223 28711 14251 28716
rect 14086 28692 14112 28695
rect 14086 28663 14112 28666
rect 14132 28148 14158 28151
rect 14132 28119 14158 28122
rect 14138 26247 14152 28119
rect 14132 26244 14158 26247
rect 14132 26215 14158 26218
rect 13994 24918 14020 24921
rect 13994 24889 14020 24892
rect 14000 24615 14014 24889
rect 13994 24612 14020 24615
rect 13994 24583 14020 24586
rect 14000 24445 14014 24583
rect 13994 24442 14020 24445
rect 13994 24413 14020 24416
rect 13994 24340 14020 24343
rect 13994 24311 14020 24314
rect 14000 24071 14014 24311
rect 13994 24068 14020 24071
rect 13994 24039 14020 24042
rect 13994 22368 14020 22371
rect 13994 22339 14020 22342
rect 14000 18563 14014 22339
rect 14086 21824 14112 21827
rect 14086 21795 14112 21798
rect 14092 20248 14106 21795
rect 14085 20244 14113 20248
rect 14085 20211 14113 20216
rect 14086 18900 14112 18903
rect 14086 18871 14112 18874
rect 14092 18631 14106 18871
rect 14086 18628 14112 18631
rect 14086 18599 14112 18602
rect 13994 18560 14020 18563
rect 14020 18540 14106 18554
rect 13994 18531 14020 18534
rect 13994 18458 14020 18461
rect 13994 18429 14020 18432
rect 13948 18084 13974 18087
rect 13948 18055 13974 18058
rect 13902 17472 13928 17475
rect 13902 17443 13928 17446
rect 13954 17305 13968 18055
rect 13948 17302 13974 17305
rect 13948 17273 13974 17276
rect 13856 16724 13882 16727
rect 13856 16695 13882 16698
rect 13586 15863 13646 15877
rect 13028 15670 13054 15673
rect 13028 15641 13054 15644
rect 13258 15364 13284 15367
rect 13258 15335 13284 15338
rect 13028 15160 13054 15163
rect 13028 15131 13054 15134
rect 13034 14925 13048 15131
rect 13028 14922 13054 14925
rect 13028 14893 13054 14896
rect 13034 13097 13048 14893
rect 13264 14536 13278 15335
rect 13396 15024 13422 15027
rect 13396 14995 13422 14998
rect 13402 14823 13416 14995
rect 13396 14820 13422 14823
rect 13396 14791 13422 14794
rect 13534 14820 13560 14823
rect 13534 14791 13560 14794
rect 13540 14653 13554 14791
rect 13534 14650 13560 14653
rect 13534 14621 13560 14624
rect 13257 14532 13285 14536
rect 13257 14499 13285 14504
rect 13264 14279 13278 14499
rect 13258 14276 13284 14279
rect 13258 14247 13284 14250
rect 13586 13191 13600 15863
rect 13672 15568 13698 15571
rect 13672 15539 13698 15542
rect 13678 14891 13692 15539
rect 13810 15364 13836 15367
rect 13810 15335 13836 15338
rect 13718 15092 13744 15095
rect 13718 15063 13744 15066
rect 13672 14888 13698 14891
rect 13672 14859 13698 14862
rect 13724 14823 13738 15063
rect 13816 14857 13830 15335
rect 13810 14854 13836 14857
rect 13810 14825 13836 14828
rect 13718 14820 13744 14823
rect 13718 14791 13744 14794
rect 13810 14786 13836 14789
rect 13810 14757 13836 14760
rect 13816 14279 13830 14757
rect 13810 14276 13836 14279
rect 13810 14247 13836 14250
rect 13580 13188 13606 13191
rect 13580 13159 13606 13162
rect 13034 13083 13094 13097
rect 12988 13015 13048 13029
rect 13034 12987 13048 13015
rect 13028 12984 13054 12987
rect 13028 12955 13054 12958
rect 12936 12950 12962 12953
rect 12936 12921 12962 12924
rect 12798 12916 12824 12919
rect 12798 12887 12824 12890
rect 12614 12576 12640 12579
rect 12614 12547 12640 12550
rect 12620 12443 12634 12547
rect 12614 12440 12640 12443
rect 12614 12411 12640 12414
rect 12804 12307 12818 12887
rect 12890 12406 12916 12409
rect 12942 12400 12956 12921
rect 13034 12647 13048 12955
rect 13028 12644 13054 12647
rect 13028 12615 13054 12618
rect 12916 12386 12956 12400
rect 12890 12377 12916 12380
rect 12798 12304 12824 12307
rect 12798 12275 12824 12278
rect 12804 12103 12818 12275
rect 12798 12100 12824 12103
rect 12798 12071 12824 12074
rect 12804 11865 12818 12071
rect 12896 12069 12910 12377
rect 12890 12066 12916 12069
rect 12890 12037 12916 12040
rect 12798 11862 12824 11865
rect 12896 11856 12910 12037
rect 13027 11948 13055 11952
rect 13027 11915 13055 11920
rect 13034 11899 13048 11915
rect 13028 11896 13054 11899
rect 13028 11867 13054 11870
rect 12936 11862 12962 11865
rect 12896 11842 12936 11856
rect 12798 11833 12824 11836
rect 12936 11833 12962 11836
rect 12804 11593 12818 11833
rect 12798 11590 12824 11593
rect 12798 11561 12824 11564
rect 12942 11525 12956 11833
rect 12982 11556 13008 11559
rect 13034 11550 13048 11867
rect 13080 11661 13094 13083
rect 13862 12428 13876 16695
rect 13954 16455 13968 17273
rect 13948 16452 13974 16455
rect 13948 16423 13974 16426
rect 13954 15367 13968 16423
rect 14000 15877 14014 18429
rect 14040 16962 14066 16965
rect 14040 16933 14066 16936
rect 14046 16829 14060 16933
rect 14040 16826 14066 16829
rect 14040 16797 14066 16800
rect 14092 16727 14106 18540
rect 14086 16724 14112 16727
rect 14086 16695 14112 16698
rect 14000 15863 14060 15877
rect 13948 15364 13974 15367
rect 13948 15335 13974 15338
rect 13954 14789 13968 15335
rect 14046 15333 14060 15863
rect 14040 15330 14066 15333
rect 14040 15301 14066 15304
rect 13948 14786 13974 14789
rect 13948 14757 13974 14760
rect 13902 14752 13928 14755
rect 13902 14723 13928 14726
rect 13908 12613 13922 14723
rect 14046 13720 14060 15301
rect 14039 13716 14067 13720
rect 14039 13683 14067 13688
rect 14138 13652 14152 26215
rect 14178 24442 14204 24445
rect 14178 24413 14204 24416
rect 14184 24071 14198 24413
rect 14178 24068 14204 24071
rect 14178 24039 14204 24042
rect 14230 23051 14244 28711
rect 14322 28185 14336 28867
rect 14362 28726 14388 28729
rect 14362 28697 14388 28700
rect 14368 28185 14382 28697
rect 14500 28386 14526 28389
rect 14500 28357 14526 28360
rect 14506 28253 14520 28357
rect 14500 28250 14526 28253
rect 14500 28221 14526 28224
rect 14316 28182 14342 28185
rect 14316 28153 14342 28156
rect 14362 28182 14388 28185
rect 14362 28153 14388 28156
rect 14454 28182 14480 28185
rect 14454 28153 14480 28156
rect 14500 28182 14526 28185
rect 14500 28153 14526 28156
rect 14546 28182 14572 28185
rect 14546 28153 14572 28156
rect 14460 27947 14474 28153
rect 14454 27944 14480 27947
rect 14454 27915 14480 27918
rect 14506 27879 14520 28153
rect 14500 27876 14526 27879
rect 14500 27847 14526 27850
rect 14552 27675 14566 28153
rect 14546 27672 14572 27675
rect 14546 27643 14572 27646
rect 14598 27301 14612 28867
rect 14914 28760 14940 28763
rect 14914 28731 14940 28734
rect 14920 28423 14934 28731
rect 15466 28454 15492 28457
rect 15466 28425 15492 28428
rect 14914 28420 14940 28423
rect 14914 28391 14940 28394
rect 15282 28250 15308 28253
rect 15282 28221 15308 28224
rect 15288 27879 15302 28221
rect 15472 28185 15486 28425
rect 15466 28182 15492 28185
rect 15466 28153 15492 28156
rect 15282 27876 15308 27879
rect 15282 27847 15308 27850
rect 15288 27641 15302 27847
rect 15702 27649 15716 29003
rect 15794 28967 15808 29241
rect 15886 29171 15900 29785
rect 16248 29712 16274 29715
rect 16248 29683 16274 29686
rect 16202 29508 16228 29511
rect 16202 29479 16228 29482
rect 15926 29236 15952 29239
rect 15926 29207 15952 29210
rect 15880 29168 15906 29171
rect 15880 29139 15906 29142
rect 15886 28967 15900 29139
rect 15788 28964 15814 28967
rect 15788 28935 15814 28938
rect 15880 28964 15906 28967
rect 15880 28935 15906 28938
rect 15742 28930 15768 28933
rect 15742 28901 15768 28904
rect 15748 28729 15762 28901
rect 15742 28726 15768 28729
rect 15742 28697 15768 28700
rect 15880 28726 15906 28729
rect 15880 28697 15906 28700
rect 15748 28457 15762 28697
rect 15742 28454 15768 28457
rect 15742 28425 15768 28428
rect 15834 28420 15860 28423
rect 15834 28391 15860 28394
rect 15840 28185 15854 28391
rect 15834 28182 15860 28185
rect 15834 28153 15860 28156
rect 15886 27675 15900 28697
rect 15932 28355 15946 29207
rect 16208 28967 16222 29479
rect 16254 28967 16268 29683
rect 16340 29542 16366 29545
rect 16340 29513 16366 29516
rect 16294 29270 16320 29273
rect 16294 29241 16320 29244
rect 16300 29069 16314 29241
rect 16294 29066 16320 29069
rect 16294 29037 16320 29040
rect 16202 28964 16228 28967
rect 16202 28935 16228 28938
rect 16248 28964 16274 28967
rect 16248 28935 16274 28938
rect 16208 28797 16222 28935
rect 16202 28794 16228 28797
rect 16202 28765 16228 28768
rect 16346 28661 16360 29513
rect 16386 29440 16412 29443
rect 16386 29411 16412 29414
rect 16392 28967 16406 29411
rect 16386 28964 16412 28967
rect 16386 28935 16412 28938
rect 17030 28964 17056 28967
rect 17030 28935 17056 28938
rect 17076 28964 17102 28967
rect 17076 28935 17102 28938
rect 17036 28797 17050 28935
rect 17030 28794 17056 28797
rect 17030 28765 17056 28768
rect 16340 28658 16366 28661
rect 16340 28629 16366 28632
rect 16846 28658 16872 28661
rect 16846 28629 16872 28632
rect 15972 28454 15998 28457
rect 15972 28425 15998 28428
rect 15926 28352 15952 28355
rect 15926 28323 15952 28326
rect 15978 28219 15992 28425
rect 16708 28420 16734 28423
rect 16708 28391 16734 28394
rect 15972 28216 15998 28219
rect 15972 28187 15998 28190
rect 16714 28185 16728 28391
rect 16852 28355 16866 28629
rect 17036 28457 17050 28765
rect 17030 28454 17056 28457
rect 17030 28425 17056 28428
rect 16846 28352 16872 28355
rect 16846 28323 16872 28326
rect 17082 28185 17096 28935
rect 17168 28930 17194 28933
rect 17168 28901 17194 28904
rect 17674 28930 17700 28933
rect 17674 28901 17700 28904
rect 17174 28491 17188 28901
rect 17214 28896 17240 28899
rect 17214 28867 17240 28870
rect 17220 28695 17234 28867
rect 17398 28726 17424 28729
rect 17398 28697 17424 28700
rect 17214 28692 17240 28695
rect 17214 28663 17240 28666
rect 17168 28488 17194 28491
rect 17168 28459 17194 28462
rect 17174 28185 17188 28459
rect 16708 28182 16734 28185
rect 16708 28153 16734 28156
rect 17076 28182 17102 28185
rect 17076 28153 17102 28156
rect 17168 28182 17194 28185
rect 17168 28153 17194 28156
rect 17220 28176 17234 28663
rect 17260 28624 17286 28627
rect 17260 28595 17286 28598
rect 17266 28423 17280 28595
rect 17260 28420 17286 28423
rect 17260 28391 17286 28394
rect 17306 28250 17332 28253
rect 17306 28221 17332 28224
rect 17260 28182 17286 28185
rect 17220 28162 17260 28176
rect 17220 27913 17234 28162
rect 17260 28153 17286 28156
rect 17214 27910 17240 27913
rect 17214 27881 17240 27884
rect 15880 27672 15906 27675
rect 15144 27638 15170 27641
rect 15144 27609 15170 27612
rect 15282 27638 15308 27641
rect 15702 27638 15854 27649
rect 15906 27646 15946 27649
rect 15880 27643 15946 27646
rect 15702 27635 15742 27638
rect 15282 27609 15308 27612
rect 15768 27635 15854 27638
rect 15886 27635 15946 27643
rect 15742 27609 15768 27612
rect 14960 27400 14986 27403
rect 14960 27371 14986 27374
rect 14592 27298 14618 27301
rect 14592 27269 14618 27272
rect 14598 27131 14612 27269
rect 14966 27131 14980 27371
rect 15052 27264 15078 27267
rect 15052 27235 15078 27238
rect 15098 27264 15124 27267
rect 15098 27235 15124 27238
rect 14592 27128 14618 27131
rect 14592 27099 14618 27102
rect 14960 27128 14986 27131
rect 14960 27099 14986 27102
rect 15006 27128 15032 27131
rect 15006 27099 15032 27102
rect 14592 27060 14618 27063
rect 14592 27031 14618 27034
rect 14598 26825 14612 27031
rect 14592 26822 14618 26825
rect 14592 26793 14618 26796
rect 14960 26516 14986 26519
rect 14960 26487 14986 26490
rect 14966 26281 14980 26487
rect 14454 26278 14480 26281
rect 14454 26249 14480 26252
rect 14960 26278 14986 26281
rect 14960 26249 14986 26252
rect 14460 26179 14474 26249
rect 14454 26176 14480 26179
rect 14454 26147 14480 26150
rect 14460 26009 14474 26147
rect 14454 26006 14480 26009
rect 14454 25977 14480 25980
rect 14408 24816 14434 24819
rect 14408 24787 14434 24790
rect 14414 24249 14428 24787
rect 14460 24343 14474 25977
rect 14914 25156 14940 25159
rect 14914 25127 14940 25130
rect 14500 25088 14526 25091
rect 14500 25059 14526 25062
rect 14506 24615 14520 25059
rect 14920 24955 14934 25127
rect 14914 24952 14940 24955
rect 14914 24923 14940 24926
rect 14776 24918 14802 24921
rect 14776 24889 14802 24892
rect 14782 24649 14796 24889
rect 14868 24816 14894 24819
rect 14868 24787 14894 24790
rect 14776 24646 14802 24649
rect 14776 24617 14802 24620
rect 14874 24615 14888 24787
rect 14920 24649 14934 24923
rect 14914 24646 14940 24649
rect 14914 24617 14940 24620
rect 14500 24612 14526 24615
rect 14500 24583 14526 24586
rect 14822 24612 14848 24615
rect 14822 24583 14848 24586
rect 14868 24612 14894 24615
rect 14868 24583 14894 24586
rect 14454 24340 14480 24343
rect 14454 24311 14480 24314
rect 14414 24235 14474 24249
rect 14224 23048 14250 23051
rect 14224 23019 14250 23022
rect 14408 22946 14434 22949
rect 14408 22917 14434 22920
rect 14362 21824 14388 21827
rect 14322 21804 14362 21818
rect 14224 21654 14250 21657
rect 14224 21625 14250 21628
rect 14178 21620 14204 21623
rect 14178 21591 14204 21594
rect 14184 21351 14198 21591
rect 14178 21348 14204 21351
rect 14178 21319 14204 21322
rect 14184 20909 14198 21319
rect 14230 21317 14244 21625
rect 14224 21314 14250 21317
rect 14224 21285 14250 21288
rect 14270 21076 14296 21079
rect 14270 21047 14296 21050
rect 14178 20906 14204 20909
rect 14178 20877 14204 20880
rect 14224 20600 14250 20603
rect 14224 20571 14250 20574
rect 14230 20365 14244 20571
rect 14224 20362 14250 20365
rect 14224 20333 14250 20336
rect 14224 20192 14250 20195
rect 14224 20163 14250 20166
rect 14230 20044 14244 20163
rect 14223 20040 14251 20044
rect 14223 20007 14251 20012
rect 14230 15877 14244 20007
rect 14276 19327 14290 21047
rect 14322 20263 14336 21804
rect 14362 21795 14388 21798
rect 14414 21317 14428 22917
rect 14408 21314 14434 21317
rect 14408 21285 14434 21288
rect 14414 21079 14428 21285
rect 14408 21076 14434 21079
rect 14408 21047 14434 21050
rect 14460 20288 14474 24235
rect 14500 24068 14526 24071
rect 14500 24039 14526 24042
rect 14506 22983 14520 24039
rect 14638 23762 14664 23765
rect 14638 23733 14664 23736
rect 14644 23357 14658 23733
rect 14638 23354 14664 23357
rect 14638 23325 14664 23328
rect 14684 23014 14710 23017
rect 14684 22985 14710 22988
rect 14500 22980 14526 22983
rect 14500 22951 14526 22954
rect 14690 22813 14704 22985
rect 14546 22810 14572 22813
rect 14546 22781 14572 22784
rect 14684 22810 14710 22813
rect 14684 22781 14710 22784
rect 14500 22436 14526 22439
rect 14500 22407 14526 22410
rect 14506 21895 14520 22407
rect 14500 21892 14526 21895
rect 14500 21863 14526 21866
rect 14552 21691 14566 22781
rect 14828 22745 14842 24583
rect 14874 24071 14888 24583
rect 14914 24408 14940 24411
rect 14914 24379 14940 24382
rect 14868 24068 14894 24071
rect 14868 24039 14894 24042
rect 14920 23289 14934 24379
rect 14966 23833 14980 26249
rect 15012 25941 15026 27099
rect 15058 26859 15072 27235
rect 15104 27063 15118 27235
rect 15150 27165 15164 27609
rect 15466 27604 15492 27607
rect 15466 27575 15492 27578
rect 15144 27162 15170 27165
rect 15144 27133 15170 27136
rect 15098 27060 15124 27063
rect 15098 27031 15124 27034
rect 15052 26856 15078 26859
rect 15052 26827 15078 26830
rect 15150 26791 15164 27133
rect 15472 27131 15486 27575
rect 15466 27128 15492 27131
rect 15466 27099 15492 27102
rect 15144 26788 15170 26791
rect 15144 26759 15170 26762
rect 15840 26587 15854 27635
rect 15834 26584 15860 26587
rect 15834 26555 15860 26558
rect 15932 26553 15946 27635
rect 16432 27332 16458 27335
rect 16432 27303 16458 27306
rect 17168 27332 17194 27335
rect 17168 27303 17194 27306
rect 16340 27094 16366 27097
rect 16340 27065 16366 27068
rect 15926 26550 15952 26553
rect 15926 26521 15952 26524
rect 15006 25938 15032 25941
rect 15006 25909 15032 25912
rect 15012 25159 15026 25909
rect 15932 25635 15946 26521
rect 16346 26519 16360 27065
rect 16340 26516 16366 26519
rect 16340 26487 16366 26490
rect 16202 26448 16228 26451
rect 16202 26419 16228 26422
rect 16340 26448 16366 26451
rect 16340 26419 16366 26422
rect 16208 26213 16222 26419
rect 16346 26349 16360 26419
rect 16340 26346 16366 26349
rect 16340 26317 16366 26320
rect 16294 26244 16320 26247
rect 16294 26215 16320 26218
rect 16202 26210 16228 26213
rect 16202 26181 16228 26184
rect 16300 25805 16314 26215
rect 16438 26179 16452 27303
rect 16478 27264 16504 27267
rect 16478 27235 16504 27238
rect 16570 27264 16596 27267
rect 16570 27235 16596 27238
rect 16484 27097 16498 27235
rect 16576 27131 16590 27235
rect 16570 27128 16596 27131
rect 16570 27099 16596 27102
rect 16478 27094 16504 27097
rect 16478 27065 16504 27068
rect 16616 26992 16642 26995
rect 16616 26963 16642 26966
rect 16622 26791 16636 26963
rect 16616 26788 16642 26791
rect 16616 26759 16642 26762
rect 17174 26723 17188 27303
rect 17312 27063 17326 28221
rect 17404 28219 17418 28697
rect 17444 28692 17470 28695
rect 17444 28663 17470 28666
rect 17582 28692 17608 28695
rect 17582 28663 17608 28666
rect 17450 28389 17464 28663
rect 17444 28386 17470 28389
rect 17444 28357 17470 28360
rect 17588 28253 17602 28663
rect 17680 28627 17694 28901
rect 18088 28794 18114 28797
rect 18088 28765 18114 28768
rect 17674 28624 17700 28627
rect 17674 28595 17700 28598
rect 17582 28250 17608 28253
rect 17582 28221 17608 28224
rect 17398 28216 17424 28219
rect 17398 28187 17424 28190
rect 17444 28114 17470 28117
rect 17444 28085 17470 28088
rect 17450 27913 17464 28085
rect 17444 27910 17470 27913
rect 17444 27881 17470 27884
rect 17680 27879 17694 28595
rect 17904 28352 17930 28355
rect 17904 28323 17930 28326
rect 17910 28151 17924 28323
rect 18094 28185 18108 28765
rect 19244 28457 19258 33000
rect 20532 29077 20546 33000
rect 20486 29063 20546 29077
rect 20158 28692 20184 28695
rect 20158 28663 20184 28666
rect 20296 28692 20322 28695
rect 20296 28663 20322 28666
rect 19238 28454 19264 28457
rect 19238 28425 19264 28428
rect 18502 28386 18528 28389
rect 18502 28357 18528 28360
rect 18088 28182 18114 28185
rect 18088 28153 18114 28156
rect 17812 28148 17838 28151
rect 17812 28119 17838 28122
rect 17904 28148 17930 28151
rect 17904 28119 17930 28122
rect 17818 27981 17832 28119
rect 17812 27978 17838 27981
rect 17812 27949 17838 27952
rect 17674 27876 17700 27879
rect 17674 27847 17700 27850
rect 17444 27808 17470 27811
rect 17444 27779 17470 27782
rect 17306 27060 17332 27063
rect 17306 27031 17332 27034
rect 17168 26720 17194 26723
rect 17168 26691 17194 26694
rect 17174 26553 17188 26691
rect 17214 26584 17240 26587
rect 17214 26555 17240 26558
rect 17168 26550 17194 26553
rect 17168 26521 17194 26524
rect 16432 26176 16458 26179
rect 16432 26147 16458 26150
rect 16294 25802 16320 25805
rect 16294 25773 16320 25776
rect 17122 25734 17148 25737
rect 17122 25705 17148 25708
rect 16708 25700 16734 25703
rect 16708 25671 16734 25674
rect 15926 25632 15952 25635
rect 15926 25603 15952 25606
rect 15052 25190 15078 25193
rect 15052 25161 15078 25164
rect 15006 25156 15032 25159
rect 15006 25127 15032 25130
rect 15012 24989 15026 25127
rect 15006 24986 15032 24989
rect 15006 24957 15032 24960
rect 15058 24887 15072 25161
rect 16156 25156 16182 25159
rect 16156 25127 16182 25130
rect 15880 24986 15906 24989
rect 15880 24957 15906 24960
rect 15886 24921 15900 24957
rect 15880 24918 15906 24921
rect 15880 24889 15906 24892
rect 15052 24884 15078 24887
rect 15052 24855 15078 24858
rect 15058 24649 15072 24855
rect 16018 24816 16044 24819
rect 16018 24787 16044 24790
rect 15052 24646 15078 24649
rect 15052 24617 15078 24620
rect 15650 24578 15676 24581
rect 15650 24549 15676 24552
rect 15052 24544 15078 24547
rect 15052 24515 15078 24518
rect 15058 23833 15072 24515
rect 15144 24374 15170 24377
rect 15144 24345 15170 24348
rect 14960 23830 14986 23833
rect 14960 23801 14986 23804
rect 15052 23830 15078 23833
rect 15052 23801 15078 23804
rect 14966 23323 14980 23801
rect 14960 23320 14986 23323
rect 14960 23291 14986 23294
rect 14914 23286 14940 23289
rect 14914 23257 14940 23260
rect 14966 22983 14980 23291
rect 15006 23252 15032 23255
rect 15006 23223 15032 23226
rect 14960 22980 14986 22983
rect 14960 22951 14986 22954
rect 14966 22813 14980 22951
rect 14960 22810 14986 22813
rect 14960 22781 14986 22784
rect 14822 22742 14848 22745
rect 14822 22713 14848 22716
rect 14960 22742 14986 22745
rect 14960 22713 14986 22716
rect 14914 22708 14940 22711
rect 14914 22679 14940 22682
rect 14776 22266 14802 22269
rect 14776 22237 14802 22240
rect 14546 21688 14572 21691
rect 14546 21659 14572 21662
rect 14460 20274 14497 20288
rect 14316 20260 14342 20263
rect 14423 20260 14449 20263
rect 14414 20248 14423 20254
rect 14316 20231 14342 20234
rect 14407 20244 14423 20248
rect 14435 20231 14449 20234
rect 14483 20237 14497 20274
rect 14483 20223 14520 20237
rect 14407 20211 14435 20216
rect 14362 20192 14388 20195
rect 14423 20192 14449 20195
rect 14362 20163 14388 20166
rect 14414 20166 14423 20186
rect 14414 20163 14449 20166
rect 14368 20093 14382 20163
rect 14362 20090 14388 20093
rect 14362 20061 14388 20064
rect 14362 19818 14388 19821
rect 14414 19812 14428 20163
rect 14388 19798 14428 19812
rect 14362 19789 14388 19792
rect 14506 19761 14520 20223
rect 14460 19747 14520 19761
rect 14276 19313 14428 19327
rect 14316 18968 14342 18971
rect 14316 18939 14342 18942
rect 14322 18631 14336 18939
rect 14316 18628 14342 18631
rect 14316 18599 14342 18602
rect 14316 17200 14342 17203
rect 14316 17171 14342 17174
rect 14270 16928 14296 16931
rect 14270 16899 14296 16902
rect 14276 16795 14290 16899
rect 14270 16792 14296 16795
rect 14270 16763 14296 16766
rect 14322 16761 14336 17171
rect 14316 16758 14342 16761
rect 14316 16729 14342 16732
rect 14230 15863 14290 15877
rect 14276 15095 14290 15863
rect 14270 15092 14296 15095
rect 14270 15063 14296 15066
rect 14178 14854 14204 14857
rect 14178 14825 14204 14828
rect 14184 14551 14198 14825
rect 14224 14786 14250 14789
rect 14224 14757 14250 14760
rect 14230 14585 14244 14757
rect 14224 14582 14250 14585
rect 14224 14553 14250 14556
rect 14178 14548 14204 14551
rect 14178 14519 14204 14522
rect 14178 13732 14204 13735
rect 14178 13703 14204 13706
rect 14131 13648 14159 13652
rect 14131 13615 14159 13620
rect 14184 13463 14198 13703
rect 14178 13460 14204 13463
rect 14178 13431 14204 13434
rect 14040 12746 14066 12749
rect 14040 12717 14066 12720
rect 13902 12610 13928 12613
rect 13902 12581 13928 12584
rect 13994 12576 14020 12579
rect 13994 12547 14020 12550
rect 13855 12424 13883 12428
rect 13855 12391 13883 12396
rect 13165 12356 13193 12360
rect 13165 12323 13193 12328
rect 13172 12069 13186 12323
rect 13862 12137 13876 12391
rect 14000 12205 14014 12547
rect 13994 12202 14020 12205
rect 13994 12173 14020 12176
rect 13856 12134 13882 12137
rect 13856 12105 13882 12108
rect 13166 12066 13192 12069
rect 13166 12037 13192 12040
rect 13172 11763 13186 12037
rect 14046 11797 14060 12717
rect 14224 12304 14250 12307
rect 14224 12275 14250 12278
rect 14276 12281 14290 15063
rect 14414 14789 14428 19313
rect 14460 18597 14474 19747
rect 14454 18594 14480 18597
rect 14454 18565 14480 18568
rect 14460 18461 14474 18565
rect 14454 18458 14480 18461
rect 14454 18429 14480 18432
rect 14454 18356 14480 18359
rect 14454 18327 14480 18330
rect 14460 18189 14474 18327
rect 14454 18186 14480 18189
rect 14454 18157 14480 18160
rect 14460 17993 14474 18157
rect 14460 17979 14520 17993
rect 14454 17472 14480 17475
rect 14454 17443 14480 17446
rect 14460 17339 14474 17443
rect 14454 17336 14480 17339
rect 14454 17307 14480 17310
rect 14506 17271 14520 17979
rect 14500 17268 14526 17271
rect 14500 17239 14526 17242
rect 14454 16758 14480 16761
rect 14552 16752 14566 21659
rect 14782 20569 14796 22237
rect 14868 20736 14894 20739
rect 14868 20707 14894 20710
rect 14874 20569 14888 20707
rect 14776 20566 14802 20569
rect 14776 20537 14802 20540
rect 14868 20566 14894 20569
rect 14868 20537 14894 20540
rect 14730 20260 14756 20263
rect 14730 20231 14756 20234
rect 14736 19787 14750 20231
rect 14730 19784 14756 19787
rect 14730 19755 14756 19758
rect 14592 18934 14618 18937
rect 14592 18905 14618 18908
rect 14598 18140 14612 18905
rect 14684 18288 14710 18291
rect 14684 18259 14710 18262
rect 14690 18189 14704 18259
rect 14684 18186 14710 18189
rect 14684 18157 14710 18160
rect 14591 18136 14619 18140
rect 14591 18103 14619 18108
rect 14684 18084 14710 18087
rect 14684 18055 14710 18058
rect 14690 17917 14704 18055
rect 14684 17914 14710 17917
rect 14684 17885 14710 17888
rect 14736 16999 14750 19755
rect 14920 18616 14934 22679
rect 14966 22201 14980 22713
rect 14960 22198 14986 22201
rect 14960 22169 14986 22172
rect 14966 21895 14980 22169
rect 14960 21892 14986 21895
rect 14960 21863 14986 21866
rect 15012 20707 15026 23223
rect 15098 23014 15124 23017
rect 15098 22985 15124 22988
rect 15052 22436 15078 22439
rect 15052 22407 15078 22410
rect 15058 22201 15072 22407
rect 15052 22198 15078 22201
rect 15052 22169 15078 22172
rect 15104 22084 15118 22985
rect 15150 22711 15164 24345
rect 15190 23796 15216 23799
rect 15190 23767 15216 23770
rect 15144 22708 15170 22711
rect 15144 22679 15170 22682
rect 15144 22266 15170 22269
rect 15144 22237 15170 22240
rect 15097 22080 15125 22084
rect 15097 22047 15125 22052
rect 15012 20693 15072 20707
rect 15006 20498 15032 20501
rect 15006 20469 15032 20472
rect 15012 20025 15026 20469
rect 15006 20022 15032 20025
rect 15006 19993 15032 19996
rect 14960 19002 14986 19005
rect 14960 18973 14986 18976
rect 14913 18612 14941 18616
rect 14913 18579 14941 18584
rect 14920 18333 14934 18579
rect 14782 18319 14934 18333
rect 14782 18087 14796 18319
rect 14868 18152 14894 18155
rect 14966 18146 14980 18973
rect 14894 18132 14980 18146
rect 14868 18123 14894 18126
rect 14776 18084 14802 18087
rect 14802 18058 14842 18061
rect 14776 18055 14842 18058
rect 14782 18047 14842 18055
rect 14730 16996 14756 16999
rect 14730 16967 14756 16970
rect 14776 16962 14802 16965
rect 14776 16933 14802 16936
rect 14454 16729 14480 16732
rect 14506 16738 14566 16752
rect 14637 16776 14665 16780
rect 14637 16743 14638 16748
rect 14460 16285 14474 16729
rect 14506 16455 14520 16738
rect 14664 16743 14665 16748
rect 14638 16729 14664 16732
rect 14545 16708 14573 16712
rect 14545 16675 14546 16680
rect 14572 16675 14573 16680
rect 14546 16661 14572 16664
rect 14500 16452 14526 16455
rect 14500 16423 14526 16426
rect 14454 16282 14480 16285
rect 14454 16253 14480 16256
rect 14506 15877 14520 16423
rect 14460 15863 14520 15877
rect 14408 14786 14434 14789
rect 14408 14757 14434 14760
rect 14362 13494 14388 13497
rect 14414 13488 14428 14757
rect 14460 14109 14474 15863
rect 14552 15148 14566 16661
rect 14782 16557 14796 16933
rect 14776 16554 14802 16557
rect 14776 16525 14802 16528
rect 14828 15877 14842 18047
rect 14868 16928 14894 16931
rect 14868 16899 14894 16902
rect 14874 16795 14888 16899
rect 14868 16792 14894 16795
rect 14868 16763 14894 16766
rect 14644 15863 14842 15877
rect 14545 15144 14573 15148
rect 14500 15126 14526 15129
rect 14545 15111 14573 15116
rect 14500 15097 14526 15100
rect 14506 14381 14520 15097
rect 14500 14378 14526 14381
rect 14500 14349 14526 14352
rect 14454 14106 14480 14109
rect 14454 14077 14480 14080
rect 14460 13701 14474 14077
rect 14592 13936 14618 13939
rect 14592 13907 14618 13910
rect 14500 13732 14526 13735
rect 14500 13703 14526 13706
rect 14545 13716 14573 13720
rect 14454 13698 14480 13701
rect 14454 13669 14480 13672
rect 14388 13474 14428 13488
rect 14454 13494 14480 13497
rect 14362 13465 14388 13468
rect 14506 13488 14520 13703
rect 14545 13683 14573 13688
rect 14552 13531 14566 13683
rect 14546 13528 14572 13531
rect 14546 13499 14572 13502
rect 14480 13474 14520 13488
rect 14454 13465 14480 13468
rect 14316 13460 14342 13463
rect 14316 13431 14342 13434
rect 14322 12375 14336 13431
rect 14500 13188 14526 13191
rect 14500 13159 14526 13162
rect 14506 13021 14520 13159
rect 14546 13120 14572 13123
rect 14546 13091 14572 13094
rect 14500 13018 14526 13021
rect 14500 12989 14526 12992
rect 14552 12647 14566 13091
rect 14598 12681 14612 13907
rect 14644 13191 14658 15863
rect 14822 15296 14848 15299
rect 14822 15267 14848 15270
rect 14828 15163 14842 15267
rect 14822 15160 14848 15163
rect 14822 15131 14848 15134
rect 14729 13580 14757 13584
rect 14729 13547 14757 13552
rect 14684 13392 14710 13395
rect 14684 13363 14710 13366
rect 14690 13259 14704 13363
rect 14684 13256 14710 13259
rect 14684 13227 14710 13230
rect 14638 13188 14664 13191
rect 14637 13172 14638 13176
rect 14664 13172 14665 13176
rect 14637 13139 14665 13144
rect 14736 12689 14750 13547
rect 14966 13312 14980 18132
rect 15012 18087 15026 19993
rect 15058 18937 15072 20693
rect 15150 20305 15164 22237
rect 15196 21472 15210 23767
rect 15236 23456 15262 23459
rect 15236 23427 15262 23430
rect 15242 23357 15256 23427
rect 15236 23354 15262 23357
rect 15236 23325 15262 23328
rect 15236 23184 15262 23187
rect 15236 23155 15262 23158
rect 15242 22371 15256 23155
rect 15236 22368 15262 22371
rect 15236 22339 15262 22342
rect 15603 22080 15631 22084
rect 15603 22047 15631 22052
rect 15512 21722 15538 21725
rect 15512 21693 15538 21696
rect 15189 21468 15217 21472
rect 15189 21435 15217 21440
rect 15104 20291 15164 20305
rect 15104 20263 15118 20291
rect 15196 20263 15210 21435
rect 15518 20637 15532 21693
rect 15512 20634 15538 20637
rect 15512 20605 15538 20608
rect 15282 20566 15308 20569
rect 15282 20537 15308 20540
rect 15374 20566 15400 20569
rect 15374 20537 15400 20540
rect 15098 20260 15124 20263
rect 15098 20231 15124 20234
rect 15190 20260 15216 20263
rect 15190 20231 15216 20234
rect 15288 20229 15302 20537
rect 15380 20365 15394 20537
rect 15374 20362 15400 20365
rect 15374 20333 15400 20336
rect 15420 20260 15446 20263
rect 15420 20231 15446 20234
rect 15282 20226 15308 20229
rect 15282 20197 15308 20200
rect 15144 20022 15170 20025
rect 15144 19993 15170 19996
rect 15052 18934 15078 18937
rect 15052 18905 15078 18908
rect 15150 18665 15164 19993
rect 15282 18900 15308 18903
rect 15282 18871 15308 18874
rect 15144 18662 15170 18665
rect 15144 18633 15170 18636
rect 15052 18628 15078 18631
rect 15052 18599 15078 18602
rect 15058 18427 15072 18599
rect 15236 18594 15262 18597
rect 15236 18565 15262 18568
rect 15052 18424 15078 18427
rect 15052 18395 15078 18398
rect 15058 18087 15072 18395
rect 15242 18393 15256 18565
rect 15236 18390 15262 18393
rect 15236 18361 15262 18364
rect 15190 18356 15216 18359
rect 15190 18327 15216 18330
rect 15196 18121 15210 18327
rect 15190 18118 15216 18121
rect 15190 18089 15216 18092
rect 15006 18084 15032 18087
rect 15006 18055 15032 18058
rect 15052 18084 15078 18087
rect 15052 18055 15078 18058
rect 15052 18016 15078 18019
rect 15052 17987 15078 17990
rect 15006 17030 15032 17033
rect 15006 17001 15032 17004
rect 15012 16829 15026 17001
rect 15058 16829 15072 17987
rect 15144 16996 15170 16999
rect 15143 16980 15144 16984
rect 15170 16980 15171 16984
rect 15143 16947 15171 16952
rect 15006 16826 15032 16829
rect 15006 16797 15032 16800
rect 15052 16826 15078 16829
rect 15052 16797 15078 16800
rect 15196 16727 15210 18089
rect 15236 17200 15262 17203
rect 15236 17171 15262 17174
rect 15242 16999 15256 17171
rect 15236 16996 15262 16999
rect 15236 16967 15262 16970
rect 15190 16724 15216 16727
rect 15190 16695 15216 16698
rect 15288 15877 15302 18871
rect 15242 15863 15302 15877
rect 15190 15636 15216 15639
rect 15190 15607 15216 15610
rect 15196 15095 15210 15607
rect 15242 15129 15256 15863
rect 15374 15704 15400 15707
rect 15374 15675 15400 15678
rect 15282 15160 15308 15163
rect 15282 15131 15308 15134
rect 15236 15126 15262 15129
rect 15236 15097 15262 15100
rect 15190 15092 15216 15095
rect 15190 15063 15216 15066
rect 15196 14551 15210 15063
rect 15190 14548 15216 14551
rect 15190 14519 15216 14522
rect 15242 14457 15256 15097
rect 15196 14443 15256 14457
rect 15144 14378 15170 14381
rect 15144 14349 15170 14352
rect 14959 13308 14987 13312
rect 14959 13275 14987 13280
rect 14822 13256 14848 13259
rect 14822 13227 14848 13230
rect 14828 13123 14842 13227
rect 14966 13191 14980 13275
rect 14960 13188 14986 13191
rect 14960 13159 14986 13162
rect 14822 13120 14848 13123
rect 14822 13091 14848 13094
rect 14822 12848 14848 12851
rect 14822 12819 14848 12822
rect 14592 12678 14618 12681
rect 14592 12649 14618 12652
rect 14644 12675 14750 12689
rect 14546 12644 14572 12647
rect 14546 12615 14572 12618
rect 14644 12485 14658 12675
rect 14684 12644 14710 12647
rect 14684 12615 14710 12618
rect 14598 12471 14658 12485
rect 14598 12443 14612 12471
rect 14592 12440 14618 12443
rect 14592 12411 14618 12414
rect 14316 12372 14342 12375
rect 14316 12343 14342 12346
rect 14230 12103 14244 12275
rect 14276 12267 14382 12281
rect 14224 12100 14250 12103
rect 14224 12071 14250 12074
rect 14368 11865 14382 12267
rect 14690 12205 14704 12615
rect 14730 12576 14756 12579
rect 14730 12547 14756 12550
rect 14684 12202 14710 12205
rect 14684 12173 14710 12176
rect 14499 12152 14527 12156
rect 14499 12119 14527 12124
rect 14408 12100 14434 12103
rect 14408 12071 14434 12074
rect 14414 11884 14428 12071
rect 14407 11880 14435 11884
rect 14316 11862 14342 11865
rect 14316 11833 14342 11836
rect 14362 11862 14388 11865
rect 14506 11865 14520 12119
rect 14407 11847 14435 11852
rect 14500 11862 14526 11865
rect 14362 11833 14388 11836
rect 14500 11833 14526 11836
rect 14040 11794 14066 11797
rect 14040 11765 14066 11768
rect 13166 11760 13192 11763
rect 13166 11731 13192 11734
rect 14322 11661 14336 11833
rect 14368 11748 14382 11833
rect 14361 11744 14389 11748
rect 14361 11711 14389 11716
rect 13074 11658 13100 11661
rect 13074 11629 13100 11632
rect 14316 11658 14342 11661
rect 14316 11629 14342 11632
rect 13008 11536 13048 11550
rect 12982 11527 13008 11530
rect 13080 11533 13094 11629
rect 13080 11525 13186 11533
rect 12936 11522 12962 11525
rect 13080 11522 13192 11525
rect 13080 11519 13166 11522
rect 12936 11493 12962 11496
rect 13166 11493 13192 11496
rect 13948 11046 13974 11049
rect 13948 11017 13974 11020
rect 12614 11012 12640 11015
rect 12614 10983 12640 10986
rect 12620 10811 12634 10983
rect 13672 10944 13698 10947
rect 13672 10915 13698 10918
rect 13856 10944 13882 10947
rect 13856 10915 13882 10918
rect 13902 10944 13928 10947
rect 13902 10915 13928 10918
rect 12430 10808 12456 10811
rect 12430 10779 12456 10782
rect 12614 10808 12640 10811
rect 12614 10779 12640 10782
rect 11878 10740 11904 10743
rect 11878 10711 11904 10714
rect 12384 10740 12410 10743
rect 12384 10711 12410 10714
rect 10682 10672 10708 10675
rect 10682 10643 10708 10646
rect 10688 10573 10702 10643
rect 9256 10570 9282 10573
rect 9256 10541 9282 10544
rect 10682 10570 10708 10573
rect 10682 10541 10708 10544
rect 8474 10502 8500 10505
rect 8474 10473 8500 10476
rect 5668 10468 5694 10471
rect 5668 10439 5694 10442
rect 7600 10468 7626 10471
rect 7600 10439 7626 10442
rect 8336 10468 8362 10471
rect 8336 10439 8362 10442
rect 7606 10301 7620 10439
rect 7600 10298 7626 10301
rect 7600 10269 7626 10272
rect 8152 10298 8178 10301
rect 8152 10269 8178 10272
rect 7508 10196 7534 10199
rect 7508 10167 7534 10170
rect 7514 10029 7528 10167
rect 7922 10128 7948 10131
rect 7922 10099 7948 10102
rect 7508 10026 7534 10029
rect 7508 9997 7534 10000
rect 7928 9961 7942 10099
rect 7922 9958 7948 9961
rect 7922 9929 7948 9932
rect 7554 9924 7580 9927
rect 7554 9895 7580 9898
rect 7600 9924 7626 9927
rect 7600 9895 7626 9898
rect 7560 9689 7574 9895
rect 7554 9686 7580 9689
rect 7554 9657 7580 9660
rect 7606 9383 7620 9895
rect 8158 9893 8172 10269
rect 7876 9890 7902 9893
rect 7876 9861 7902 9864
rect 8152 9890 8178 9893
rect 8152 9861 8178 9864
rect 7882 9723 7896 9861
rect 7876 9720 7902 9723
rect 7876 9691 7902 9694
rect 8106 9720 8132 9723
rect 8106 9691 8132 9694
rect 7882 9655 7896 9691
rect 7876 9652 7902 9655
rect 7876 9623 7902 9626
rect 7784 9584 7810 9587
rect 7784 9555 7810 9558
rect 7790 9417 7804 9555
rect 7784 9414 7810 9417
rect 7784 9385 7810 9388
rect 7600 9380 7626 9383
rect 7600 9351 7626 9354
rect 5990 8870 6016 8873
rect 5990 8841 6016 8844
rect 6036 8870 6062 8873
rect 6036 8841 6062 8844
rect 5622 8836 5648 8839
rect 5622 8807 5648 8810
rect 5996 8057 6010 8841
rect 6042 8329 6056 8841
rect 6082 8836 6108 8839
rect 6082 8807 6108 8810
rect 6088 8329 6102 8807
rect 6358 8564 6384 8567
rect 6358 8535 6384 8538
rect 6542 8564 6568 8567
rect 6542 8535 6568 8538
rect 6036 8326 6062 8329
rect 6036 8297 6062 8300
rect 6082 8326 6108 8329
rect 6082 8297 6108 8300
rect 6082 8258 6108 8261
rect 6082 8229 6108 8232
rect 5990 8054 6016 8057
rect 5990 8025 6016 8028
rect 5996 7547 6010 8025
rect 6088 7589 6102 8229
rect 6364 8227 6378 8535
rect 6358 8224 6384 8227
rect 6358 8195 6384 8198
rect 6548 7853 6562 8535
rect 7606 8295 7620 9351
rect 7738 9346 7764 9349
rect 7738 9317 7764 9320
rect 7692 8870 7718 8873
rect 7692 8841 7718 8844
rect 7646 8768 7672 8771
rect 7646 8739 7672 8742
rect 7652 8669 7666 8739
rect 7646 8666 7672 8669
rect 7646 8637 7672 8640
rect 7698 8567 7712 8841
rect 7744 8601 7758 9317
rect 8112 8839 8126 9691
rect 8158 9349 8172 9861
rect 8342 9723 8356 10439
rect 8382 10400 8408 10403
rect 8382 10371 8408 10374
rect 8388 10233 8402 10371
rect 8382 10230 8408 10233
rect 8382 10201 8408 10204
rect 8388 9969 8402 10201
rect 8388 9961 8448 9969
rect 8388 9958 8454 9961
rect 8388 9955 8428 9958
rect 8428 9929 8454 9932
rect 8336 9720 8362 9723
rect 8336 9691 8362 9694
rect 8480 9655 8494 10473
rect 9026 10434 9052 10437
rect 9026 10405 9052 10408
rect 8934 10400 8960 10403
rect 8934 10371 8960 10374
rect 8940 10233 8954 10371
rect 9032 10267 9046 10405
rect 9262 10403 9276 10541
rect 9532 10502 9558 10505
rect 9532 10473 9558 10476
rect 9256 10400 9282 10403
rect 9256 10371 9282 10374
rect 9026 10264 9052 10267
rect 9026 10235 9052 10238
rect 8842 10230 8868 10233
rect 8842 10201 8868 10204
rect 8934 10230 8960 10233
rect 8934 10201 8960 10204
rect 8474 9652 8500 9655
rect 8474 9623 8500 9626
rect 8848 9621 8862 10201
rect 8888 9958 8914 9961
rect 8888 9929 8914 9932
rect 8894 9757 8908 9929
rect 9262 9927 9276 10371
rect 9538 10233 9552 10473
rect 9578 10434 9604 10437
rect 9578 10405 9604 10408
rect 9584 10301 9598 10405
rect 9578 10298 9604 10301
rect 9578 10269 9604 10272
rect 10544 10264 10570 10267
rect 10544 10235 10570 10238
rect 9532 10230 9558 10233
rect 9532 10201 9558 10204
rect 9538 9995 9552 10201
rect 9670 10196 9696 10199
rect 9670 10167 9696 10170
rect 9716 10196 9742 10199
rect 9716 10167 9742 10170
rect 9676 10029 9690 10167
rect 9670 10026 9696 10029
rect 9670 9997 9696 10000
rect 9532 9992 9558 9995
rect 9532 9963 9558 9966
rect 8980 9924 9006 9927
rect 8980 9895 9006 9898
rect 9256 9924 9282 9927
rect 9256 9895 9282 9898
rect 8888 9754 8914 9757
rect 8888 9725 8914 9728
rect 8934 9720 8960 9723
rect 8986 9697 9000 9895
rect 9072 9856 9098 9859
rect 9072 9827 9098 9830
rect 8960 9694 9000 9697
rect 8934 9691 9000 9694
rect 8940 9683 9000 9691
rect 8888 9652 8914 9655
rect 8888 9623 8914 9626
rect 8842 9618 8868 9621
rect 8842 9589 8868 9592
rect 8894 9417 8908 9623
rect 8888 9414 8914 9417
rect 8888 9385 8914 9388
rect 8152 9346 8178 9349
rect 8152 9317 8178 9320
rect 7876 8836 7902 8839
rect 7876 8807 7902 8810
rect 8106 8836 8132 8839
rect 8106 8807 8132 8810
rect 7830 8802 7856 8805
rect 7830 8773 7856 8776
rect 7784 8768 7810 8771
rect 7784 8739 7810 8742
rect 7738 8598 7764 8601
rect 7738 8569 7764 8572
rect 7692 8564 7718 8567
rect 7692 8535 7718 8538
rect 7600 8292 7626 8295
rect 7600 8263 7626 8266
rect 6864 8224 6890 8227
rect 6864 8195 6890 8198
rect 6588 8054 6614 8057
rect 6588 8025 6614 8028
rect 6542 7850 6568 7853
rect 6542 7821 6568 7824
rect 6594 7785 6608 8025
rect 6870 8023 6884 8195
rect 6864 8020 6890 8023
rect 6864 7991 6890 7994
rect 6818 7952 6844 7955
rect 6818 7923 6844 7926
rect 6588 7782 6614 7785
rect 6588 7753 6614 7756
rect 6824 7751 6838 7923
rect 6818 7748 6844 7751
rect 6818 7719 6844 7722
rect 6042 7575 6102 7589
rect 6174 7578 6200 7581
rect 5990 7544 6016 7547
rect 5990 7515 6016 7518
rect 5530 7204 5556 7207
rect 5530 7175 5556 7178
rect 5536 6221 5550 7175
rect 6042 7173 6056 7575
rect 6174 7549 6200 7552
rect 6082 7544 6108 7547
rect 6082 7515 6108 7518
rect 5668 7170 5694 7173
rect 5668 7141 5694 7144
rect 5944 7170 5970 7173
rect 5944 7141 5970 7144
rect 6036 7170 6062 7173
rect 6036 7141 6062 7144
rect 5674 7037 5688 7141
rect 5668 7034 5694 7037
rect 5668 7005 5694 7008
rect 5950 6357 5964 7141
rect 6088 6731 6102 7515
rect 6128 7408 6154 7411
rect 6128 7379 6154 7382
rect 6134 6969 6148 7379
rect 6180 7241 6194 7549
rect 6220 7510 6246 7513
rect 6220 7481 6246 7484
rect 6174 7238 6200 7241
rect 6174 7209 6200 7212
rect 6128 6966 6154 6969
rect 6128 6937 6154 6940
rect 6180 6909 6194 7209
rect 6134 6901 6194 6909
rect 6128 6898 6194 6901
rect 6154 6895 6194 6898
rect 6128 6869 6154 6872
rect 6082 6728 6108 6731
rect 6082 6699 6108 6702
rect 5990 6592 6016 6595
rect 5990 6563 6016 6566
rect 5944 6354 5970 6357
rect 5944 6325 5970 6328
rect 5530 6218 5556 6221
rect 5530 6189 5556 6192
rect 5950 6085 5964 6325
rect 5996 6323 6010 6563
rect 6088 6391 6102 6699
rect 6134 6595 6148 6869
rect 6226 6867 6240 7481
rect 6870 7411 6884 7991
rect 7139 7596 7167 7600
rect 7139 7563 7167 7568
rect 7146 7547 7160 7563
rect 7140 7544 7166 7547
rect 7140 7515 7166 7518
rect 7606 7411 7620 8263
rect 7698 8125 7712 8535
rect 7790 8329 7804 8739
rect 7836 8635 7850 8773
rect 7830 8632 7856 8635
rect 7830 8603 7856 8606
rect 7784 8326 7810 8329
rect 7784 8297 7810 8300
rect 7692 8122 7718 8125
rect 7692 8093 7718 8096
rect 7698 8023 7712 8093
rect 7836 8091 7850 8603
rect 7882 8601 7896 8807
rect 7922 8666 7948 8669
rect 7922 8637 7948 8640
rect 7876 8598 7902 8601
rect 7876 8569 7902 8572
rect 7876 8530 7902 8533
rect 7876 8501 7902 8504
rect 7882 8227 7896 8501
rect 7876 8224 7902 8227
rect 7876 8195 7902 8198
rect 7882 8125 7896 8195
rect 7876 8122 7902 8125
rect 7876 8093 7902 8096
rect 7738 8088 7764 8091
rect 7738 8059 7764 8062
rect 7830 8088 7856 8091
rect 7830 8059 7856 8062
rect 7646 8020 7672 8023
rect 7646 7991 7672 7994
rect 7692 8020 7718 8023
rect 7692 7991 7718 7994
rect 7652 7819 7666 7991
rect 7692 7952 7718 7955
rect 7692 7923 7718 7926
rect 7646 7816 7672 7819
rect 7646 7787 7672 7790
rect 7698 7751 7712 7923
rect 7692 7748 7718 7751
rect 7692 7719 7718 7722
rect 7698 7547 7712 7719
rect 7692 7544 7718 7547
rect 7692 7515 7718 7518
rect 7646 7510 7672 7513
rect 7646 7481 7672 7484
rect 6588 7408 6614 7411
rect 6588 7379 6614 7382
rect 6864 7408 6890 7411
rect 6864 7379 6890 7382
rect 7600 7408 7626 7411
rect 7600 7379 7626 7382
rect 6220 6864 6246 6867
rect 6220 6835 6246 6838
rect 6226 6705 6240 6835
rect 6180 6697 6240 6705
rect 6180 6694 6246 6697
rect 6180 6691 6220 6694
rect 6128 6592 6154 6595
rect 6128 6563 6154 6566
rect 6134 6493 6148 6563
rect 6128 6490 6154 6493
rect 6128 6461 6154 6464
rect 6082 6388 6108 6391
rect 6082 6359 6108 6362
rect 5990 6320 6016 6323
rect 5990 6291 6016 6294
rect 6134 6187 6148 6461
rect 6180 6425 6194 6691
rect 6220 6665 6246 6668
rect 6220 6626 6246 6629
rect 6220 6597 6246 6600
rect 6226 6459 6240 6597
rect 6220 6456 6246 6459
rect 6220 6427 6246 6430
rect 6496 6456 6522 6459
rect 6496 6427 6522 6430
rect 6174 6422 6200 6425
rect 6174 6393 6200 6396
rect 6266 6320 6292 6323
rect 6266 6291 6292 6294
rect 6128 6184 6154 6187
rect 6128 6155 6154 6158
rect 6272 6153 6286 6291
rect 6266 6150 6292 6153
rect 6266 6121 6292 6124
rect 6502 6085 6516 6427
rect 6594 6391 6608 7379
rect 7606 7241 7620 7379
rect 7600 7238 7626 7241
rect 7600 7209 7626 7212
rect 7600 7170 7626 7173
rect 7600 7141 7626 7144
rect 6772 6864 6798 6867
rect 6772 6835 6798 6838
rect 6726 6592 6752 6595
rect 6726 6563 6752 6566
rect 6732 6459 6746 6563
rect 6726 6456 6752 6459
rect 6726 6427 6752 6430
rect 6588 6388 6614 6391
rect 6588 6359 6614 6362
rect 6594 6221 6608 6359
rect 6588 6218 6614 6221
rect 6588 6189 6614 6192
rect 6778 6187 6792 6835
rect 6910 6626 6936 6629
rect 6910 6597 6936 6600
rect 6916 6221 6930 6597
rect 7606 6459 7620 7141
rect 7600 6456 7626 6459
rect 7600 6427 7626 6430
rect 7600 6388 7626 6391
rect 7600 6359 7626 6362
rect 6910 6218 6936 6221
rect 6910 6189 6936 6192
rect 6772 6184 6798 6187
rect 6772 6155 6798 6158
rect 7606 6153 7620 6359
rect 7652 6187 7666 7481
rect 7744 7453 7758 8059
rect 7836 7793 7850 8059
rect 7928 8023 7942 8637
rect 8112 8635 8126 8807
rect 8106 8632 8132 8635
rect 8106 8603 8132 8606
rect 8842 8632 8868 8635
rect 8842 8603 8868 8606
rect 8520 8598 8546 8601
rect 8520 8569 8546 8572
rect 8526 8397 8540 8569
rect 8520 8394 8546 8397
rect 8520 8365 8546 8368
rect 8848 8287 8862 8603
rect 8894 8533 8908 9385
rect 8888 8530 8914 8533
rect 8888 8501 8914 8504
rect 8980 8496 9006 8499
rect 8980 8467 9006 8470
rect 8802 8273 8862 8287
rect 8750 8258 8776 8261
rect 8750 8229 8776 8232
rect 8198 8054 8224 8057
rect 8198 8025 8224 8028
rect 7922 8020 7948 8023
rect 7922 7991 7948 7994
rect 7790 7785 7850 7793
rect 7784 7782 7850 7785
rect 7810 7779 7850 7782
rect 7784 7753 7810 7756
rect 7698 7439 7758 7453
rect 7698 7173 7712 7439
rect 7738 7408 7764 7411
rect 7738 7379 7764 7382
rect 7744 7241 7758 7379
rect 7738 7238 7764 7241
rect 7738 7209 7764 7212
rect 7692 7170 7718 7173
rect 7692 7141 7718 7144
rect 7790 6663 7804 7753
rect 7928 7717 7942 7991
rect 8204 7989 8218 8025
rect 8198 7986 8224 7989
rect 8198 7957 8224 7960
rect 8106 7952 8132 7955
rect 8106 7923 8132 7926
rect 8112 7853 8126 7923
rect 8106 7850 8132 7853
rect 8106 7821 8132 7824
rect 7922 7714 7948 7717
rect 7922 7685 7948 7688
rect 7830 7680 7856 7683
rect 7830 7651 7856 7654
rect 7784 6660 7810 6663
rect 7784 6631 7810 6634
rect 7646 6184 7672 6187
rect 7646 6155 7672 6158
rect 7600 6150 7626 6153
rect 7600 6121 7626 6124
rect 7652 6085 7666 6155
rect 7790 6119 7804 6631
rect 7784 6116 7810 6119
rect 7784 6087 7810 6090
rect 5944 6082 5970 6085
rect 5944 6053 5970 6056
rect 6496 6082 6522 6085
rect 6496 6053 6522 6056
rect 7646 6082 7672 6085
rect 7646 6053 7672 6056
rect 7508 6048 7534 6051
rect 7508 6019 7534 6022
rect 7514 5949 7528 6019
rect 7508 5946 7534 5949
rect 7508 5917 7534 5920
rect 7836 5915 7850 7651
rect 7830 5912 7856 5915
rect 7830 5883 7856 5886
rect 7738 5878 7764 5881
rect 7738 5849 7764 5852
rect 5207 5624 5235 5628
rect 5207 5591 5235 5596
rect 7744 5541 7758 5849
rect 7876 5776 7902 5779
rect 7876 5747 7902 5750
rect 7882 5609 7896 5747
rect 7876 5606 7902 5609
rect 7876 5577 7902 5580
rect 7928 5575 7942 7685
rect 8204 7683 8218 7957
rect 8756 7683 8770 8229
rect 8198 7680 8224 7683
rect 8750 7680 8776 7683
rect 8198 7651 8224 7654
rect 8749 7664 8750 7668
rect 8776 7664 8777 7668
rect 8749 7631 8777 7636
rect 8198 7442 8224 7445
rect 8198 7413 8224 7416
rect 8106 7238 8132 7241
rect 8106 7209 8132 7212
rect 8112 6969 8126 7209
rect 8106 6966 8132 6969
rect 8106 6937 8132 6940
rect 8014 6150 8040 6153
rect 8014 6121 8040 6124
rect 8020 5575 8034 6121
rect 8112 5847 8126 6937
rect 8204 6901 8218 7413
rect 8802 7309 8816 8273
rect 8842 8224 8868 8227
rect 8842 8195 8868 8198
rect 8848 7600 8862 8195
rect 8841 7596 8869 7600
rect 8841 7563 8869 7568
rect 8796 7306 8822 7309
rect 8796 7277 8822 7280
rect 8802 7037 8816 7277
rect 8888 7170 8914 7173
rect 8888 7141 8914 7144
rect 8796 7034 8822 7037
rect 8796 7005 8822 7008
rect 8894 6969 8908 7141
rect 8888 6966 8914 6969
rect 8888 6937 8914 6940
rect 8198 6898 8224 6901
rect 8198 6869 8224 6872
rect 8244 5912 8270 5915
rect 8244 5883 8270 5886
rect 8106 5844 8132 5847
rect 8106 5815 8132 5818
rect 7830 5572 7856 5575
rect 7830 5543 7856 5546
rect 7922 5572 7948 5575
rect 7922 5543 7948 5546
rect 8014 5572 8040 5575
rect 8014 5543 8040 5546
rect 7738 5538 7764 5541
rect 7738 5509 7764 5512
rect 7744 5371 7758 5509
rect 7738 5368 7764 5371
rect 7738 5339 7764 5342
rect 5529 660 5557 664
rect 5529 627 5557 632
rect 5536 0 5550 627
rect 7744 0 7758 5339
rect 7836 5031 7850 5543
rect 7928 5337 7942 5543
rect 8020 5405 8034 5543
rect 8014 5402 8040 5405
rect 8014 5373 8040 5376
rect 8250 5345 8264 5883
rect 8986 5575 9000 8467
rect 9078 8287 9092 9827
rect 9538 8873 9552 9963
rect 9578 9958 9604 9961
rect 9578 9929 9604 9932
rect 9584 9689 9598 9929
rect 9722 9927 9736 10167
rect 9716 9924 9742 9927
rect 9716 9895 9742 9898
rect 9722 9723 9736 9895
rect 10550 9893 10564 10235
rect 10314 9890 10340 9893
rect 10314 9861 10340 9864
rect 10544 9890 10570 9893
rect 10544 9861 10570 9864
rect 10820 9890 10846 9893
rect 10820 9861 10846 9864
rect 9992 9856 10018 9859
rect 9992 9827 10018 9830
rect 9716 9720 9742 9723
rect 9716 9691 9742 9694
rect 9998 9689 10012 9827
rect 9578 9686 9604 9689
rect 9578 9657 9604 9660
rect 9992 9686 10018 9689
rect 9992 9657 10018 9660
rect 10320 9655 10334 9861
rect 10314 9652 10340 9655
rect 10314 9623 10340 9626
rect 9532 8870 9558 8873
rect 9532 8841 9558 8844
rect 10360 8870 10386 8873
rect 10360 8841 10386 8844
rect 9538 8669 9552 8841
rect 9532 8666 9558 8669
rect 9532 8637 9558 8640
rect 9486 8598 9512 8601
rect 9486 8569 9512 8572
rect 9118 8564 9144 8567
rect 9118 8535 9144 8538
rect 9032 8273 9092 8287
rect 9032 7241 9046 8273
rect 9072 7510 9098 7513
rect 9072 7481 9098 7484
rect 9078 7309 9092 7481
rect 9124 7445 9138 8535
rect 9492 8397 9506 8569
rect 9486 8394 9512 8397
rect 9486 8365 9512 8368
rect 9538 8295 9552 8637
rect 9532 8292 9558 8295
rect 9532 8263 9558 8266
rect 10366 7785 10380 8841
rect 10826 8805 10840 9861
rect 11096 8870 11122 8873
rect 11096 8841 11122 8844
rect 11102 8813 11116 8841
rect 10636 8802 10662 8805
rect 10636 8773 10662 8776
rect 10820 8802 10846 8805
rect 10820 8773 10846 8776
rect 11004 8802 11030 8805
rect 11004 8773 11030 8776
rect 11056 8799 11116 8813
rect 10642 8635 10656 8773
rect 10636 8632 10662 8635
rect 10636 8603 10662 8606
rect 10452 8598 10478 8601
rect 10452 8569 10478 8572
rect 10458 8057 10472 8569
rect 10636 8564 10662 8567
rect 10636 8535 10662 8538
rect 10452 8054 10478 8057
rect 10452 8025 10478 8028
rect 10590 8054 10616 8057
rect 10590 8025 10616 8028
rect 10406 8020 10432 8023
rect 10406 7991 10432 7994
rect 10360 7782 10386 7785
rect 10360 7753 10386 7756
rect 9256 7510 9282 7513
rect 9256 7481 9282 7484
rect 9440 7510 9466 7513
rect 9440 7481 9466 7484
rect 9578 7510 9604 7513
rect 9578 7481 9604 7484
rect 9118 7442 9144 7445
rect 9118 7413 9144 7416
rect 9072 7306 9098 7309
rect 9072 7277 9098 7280
rect 9026 7238 9052 7241
rect 9026 7209 9052 7212
rect 9262 6051 9276 7481
rect 9446 7173 9460 7481
rect 9584 7207 9598 7481
rect 10366 7241 10380 7753
rect 10412 7751 10426 7991
rect 10406 7748 10432 7751
rect 10406 7719 10432 7722
rect 10412 7513 10426 7719
rect 10406 7510 10432 7513
rect 10406 7481 10432 7484
rect 10412 7453 10426 7481
rect 10412 7439 10472 7453
rect 10596 7445 10610 8025
rect 10642 8023 10656 8535
rect 10636 8020 10662 8023
rect 10636 7991 10662 7994
rect 10682 7952 10708 7955
rect 10682 7923 10708 7926
rect 10688 7785 10702 7923
rect 10682 7782 10708 7785
rect 10682 7753 10708 7756
rect 11010 7717 11024 8773
rect 11056 8601 11070 8799
rect 11050 8598 11076 8601
rect 11050 8569 11076 8572
rect 11004 7714 11030 7717
rect 11004 7685 11030 7688
rect 10406 7408 10432 7411
rect 10406 7379 10432 7382
rect 10412 7309 10426 7379
rect 10406 7306 10432 7309
rect 10406 7277 10432 7280
rect 10360 7238 10386 7241
rect 10360 7209 10386 7212
rect 9578 7204 9604 7207
rect 9578 7175 9604 7178
rect 9440 7170 9466 7173
rect 9440 7141 9466 7144
rect 9302 7136 9328 7139
rect 9302 7107 9328 7110
rect 9256 6048 9282 6051
rect 9256 6019 9282 6022
rect 9262 5915 9276 6019
rect 9256 5912 9282 5915
rect 9256 5883 9282 5886
rect 9308 5881 9322 7107
rect 9446 5881 9460 7141
rect 10458 7003 10472 7439
rect 10590 7442 10616 7445
rect 10590 7413 10616 7416
rect 10596 7275 10610 7413
rect 10728 7408 10754 7411
rect 10728 7379 10754 7382
rect 10590 7272 10616 7275
rect 10590 7243 10616 7246
rect 10734 7037 10748 7379
rect 10820 7238 10846 7241
rect 10820 7209 10846 7212
rect 10728 7034 10754 7037
rect 10728 7005 10754 7008
rect 10452 7000 10478 7003
rect 10452 6971 10478 6974
rect 10458 5915 10472 6971
rect 10826 6697 10840 7209
rect 11010 7173 11024 7685
rect 11004 7170 11030 7173
rect 11004 7141 11030 7144
rect 10820 6694 10846 6697
rect 10820 6665 10846 6668
rect 11010 6629 11024 7141
rect 11004 6626 11030 6629
rect 11004 6597 11030 6600
rect 11056 6119 11070 8569
rect 11096 8496 11122 8499
rect 11096 8467 11122 8470
rect 11102 7513 11116 8467
rect 11556 7986 11582 7989
rect 11556 7957 11582 7960
rect 11510 7714 11536 7717
rect 11510 7685 11536 7688
rect 11516 7513 11530 7685
rect 11096 7510 11122 7513
rect 11096 7481 11122 7484
rect 11510 7510 11536 7513
rect 11510 7481 11536 7484
rect 11050 6116 11076 6119
rect 11050 6087 11076 6090
rect 11102 5949 11116 7481
rect 11562 7445 11576 7957
rect 11648 7544 11674 7547
rect 11648 7515 11674 7518
rect 11556 7442 11582 7445
rect 11556 7413 11582 7416
rect 11654 7241 11668 7515
rect 11832 7510 11858 7513
rect 11832 7481 11858 7484
rect 11838 7275 11852 7481
rect 11832 7272 11858 7275
rect 11832 7243 11858 7246
rect 11648 7238 11674 7241
rect 11648 7209 11674 7212
rect 11510 7204 11536 7207
rect 11510 7175 11536 7178
rect 11142 7136 11168 7139
rect 11142 7107 11168 7110
rect 11148 6697 11162 7107
rect 11516 6901 11530 7175
rect 11838 6969 11852 7243
rect 11832 6966 11858 6969
rect 11832 6937 11858 6940
rect 11510 6898 11536 6901
rect 11510 6869 11536 6872
rect 11142 6694 11168 6697
rect 11142 6665 11168 6668
rect 11838 6629 11852 6937
rect 11832 6626 11858 6629
rect 11832 6597 11858 6600
rect 11556 6048 11582 6051
rect 11556 6019 11582 6022
rect 11096 5946 11122 5949
rect 11096 5917 11122 5920
rect 9486 5912 9512 5915
rect 9486 5883 9512 5886
rect 10452 5912 10478 5915
rect 10452 5883 10478 5886
rect 9302 5878 9328 5881
rect 9302 5849 9328 5852
rect 9440 5878 9466 5881
rect 9440 5849 9466 5852
rect 9026 5776 9052 5779
rect 9026 5747 9052 5750
rect 9032 5575 9046 5747
rect 8612 5572 8638 5575
rect 8612 5543 8638 5546
rect 8980 5572 9006 5575
rect 8980 5543 9006 5546
rect 9026 5572 9052 5575
rect 9026 5543 9052 5546
rect 8250 5337 8310 5345
rect 7922 5334 7948 5337
rect 8250 5334 8316 5337
rect 8250 5331 8290 5334
rect 7922 5305 7948 5308
rect 8290 5305 8316 5308
rect 8244 5300 8270 5303
rect 8244 5271 8270 5274
rect 8250 5031 8264 5271
rect 8618 5235 8632 5543
rect 9446 5541 9460 5849
rect 9492 5609 9506 5883
rect 11562 5881 11576 6019
rect 11838 5915 11852 6597
rect 11832 5912 11858 5915
rect 11832 5883 11858 5886
rect 9532 5878 9558 5881
rect 9532 5849 9558 5852
rect 10130 5878 10156 5881
rect 10130 5849 10156 5852
rect 10176 5878 10202 5881
rect 10176 5849 10202 5852
rect 11556 5878 11582 5881
rect 11556 5849 11582 5852
rect 9486 5606 9512 5609
rect 9486 5577 9512 5580
rect 9440 5538 9466 5541
rect 9440 5509 9466 5512
rect 9446 5337 9460 5509
rect 9538 5405 9552 5849
rect 10136 5677 10150 5849
rect 10130 5674 10156 5677
rect 10130 5645 10156 5648
rect 10182 5507 10196 5849
rect 11004 5844 11030 5847
rect 11004 5815 11030 5818
rect 10222 5572 10248 5575
rect 10222 5543 10248 5546
rect 10176 5504 10202 5507
rect 10176 5475 10202 5478
rect 9532 5402 9558 5405
rect 9532 5373 9558 5376
rect 9440 5334 9466 5337
rect 9440 5305 9466 5308
rect 10228 5269 10242 5543
rect 11010 5405 11024 5815
rect 11648 5776 11674 5779
rect 11648 5747 11674 5750
rect 11654 5609 11668 5747
rect 11648 5606 11674 5609
rect 11648 5577 11674 5580
rect 11004 5402 11030 5405
rect 11004 5373 11030 5376
rect 10222 5266 10248 5269
rect 10222 5237 10248 5240
rect 8290 5232 8316 5235
rect 8290 5203 8316 5206
rect 8612 5232 8638 5235
rect 8612 5203 8638 5206
rect 8296 5133 8310 5203
rect 8290 5130 8316 5133
rect 8290 5101 8316 5104
rect 7830 5028 7856 5031
rect 7830 4999 7856 5002
rect 8244 5028 8270 5031
rect 8244 4999 8270 5002
rect 7836 0 7850 4999
rect 11884 0 11898 10711
rect 12390 10471 12404 10711
rect 13678 10505 13692 10915
rect 13862 10505 13876 10915
rect 13908 10845 13922 10915
rect 13902 10842 13928 10845
rect 13902 10813 13928 10816
rect 13954 10573 13968 11017
rect 14500 11012 14526 11015
rect 14500 10983 14526 10986
rect 14506 10811 14520 10983
rect 14500 10808 14526 10811
rect 14500 10779 14526 10782
rect 14736 10777 14750 12547
rect 14828 12477 14842 12819
rect 14822 12474 14848 12477
rect 14822 12445 14848 12448
rect 14828 12103 14842 12445
rect 14914 12304 14940 12307
rect 14914 12275 14940 12278
rect 14920 12103 14934 12275
rect 14822 12100 14848 12103
rect 14822 12071 14848 12074
rect 14914 12100 14940 12103
rect 14914 12071 14940 12074
rect 15150 10777 15164 14349
rect 15196 14007 15210 14443
rect 15190 14004 15216 14007
rect 15190 13975 15216 13978
rect 15288 12360 15302 15131
rect 15328 14038 15354 14041
rect 15328 14009 15354 14012
rect 15334 13565 15348 14009
rect 15380 13584 15394 15675
rect 15426 14619 15440 20231
rect 15610 20059 15624 22047
rect 15604 20056 15630 20059
rect 15604 20027 15630 20030
rect 15512 18390 15538 18393
rect 15512 18361 15538 18364
rect 15466 16996 15492 16999
rect 15466 16967 15492 16970
rect 15472 16727 15486 16967
rect 15518 16837 15532 18361
rect 15557 16844 15585 16848
rect 15518 16823 15557 16837
rect 15557 16811 15585 16816
rect 15564 16795 15578 16811
rect 15558 16792 15584 16795
rect 15511 16776 15539 16780
rect 15558 16763 15584 16766
rect 15511 16743 15512 16748
rect 15538 16743 15539 16748
rect 15512 16729 15538 16732
rect 15466 16724 15492 16727
rect 15466 16695 15492 16698
rect 15472 16489 15486 16695
rect 15466 16486 15492 16489
rect 15466 16457 15492 16460
rect 15466 15670 15492 15673
rect 15466 15641 15492 15644
rect 15472 15120 15486 15641
rect 15610 15163 15624 20027
rect 15656 18903 15670 24549
rect 16024 24411 16038 24787
rect 16162 24445 16176 25127
rect 16714 24615 16728 25671
rect 17076 25190 17102 25193
rect 17076 25161 17102 25164
rect 17082 24921 17096 25161
rect 17076 24918 17102 24921
rect 17076 24889 17102 24892
rect 17082 24615 17096 24889
rect 17128 24819 17142 25705
rect 17174 25125 17188 26521
rect 17220 25703 17234 26555
rect 17259 26432 17287 26436
rect 17259 26399 17287 26404
rect 17266 26315 17280 26399
rect 17260 26312 17286 26315
rect 17260 26283 17286 26286
rect 17312 26247 17326 27031
rect 17398 26618 17424 26621
rect 17398 26589 17424 26592
rect 17306 26244 17332 26247
rect 17306 26215 17332 26218
rect 17214 25700 17240 25703
rect 17214 25671 17240 25674
rect 17260 25666 17286 25669
rect 17260 25637 17286 25640
rect 17168 25122 17194 25125
rect 17168 25093 17194 25096
rect 17174 24887 17188 25093
rect 17266 24921 17280 25637
rect 17404 25261 17418 26589
rect 17398 25258 17424 25261
rect 17398 25229 17424 25232
rect 17260 24918 17286 24921
rect 17260 24889 17286 24892
rect 17168 24884 17194 24887
rect 17168 24855 17194 24858
rect 17122 24816 17148 24819
rect 17122 24787 17148 24790
rect 16708 24612 16734 24615
rect 16708 24583 16734 24586
rect 17076 24612 17102 24615
rect 17076 24583 17102 24586
rect 16156 24442 16182 24445
rect 16156 24413 16182 24416
rect 16018 24408 16044 24411
rect 16018 24379 16044 24382
rect 16162 24377 16176 24413
rect 16156 24374 16182 24377
rect 16156 24345 16182 24348
rect 16340 24306 16366 24309
rect 16340 24277 16366 24280
rect 16294 24102 16320 24105
rect 16294 24073 16320 24076
rect 15834 23456 15860 23459
rect 15834 23427 15860 23430
rect 15696 22368 15722 22371
rect 15696 22339 15722 22342
rect 15702 18937 15716 22339
rect 15840 21657 15854 23427
rect 16300 23289 16314 24073
rect 16346 24071 16360 24277
rect 16714 24071 16728 24583
rect 16340 24068 16366 24071
rect 16340 24039 16366 24042
rect 16708 24068 16734 24071
rect 16708 24039 16734 24042
rect 16386 24000 16412 24003
rect 16386 23971 16412 23974
rect 16294 23286 16320 23289
rect 16294 23257 16320 23260
rect 16156 23218 16182 23221
rect 16156 23189 16182 23192
rect 16162 22915 16176 23189
rect 16248 22980 16274 22983
rect 16248 22951 16274 22954
rect 16156 22912 16182 22915
rect 16156 22883 16182 22886
rect 16162 21657 16176 22883
rect 16254 22745 16268 22951
rect 16248 22742 16274 22745
rect 16248 22713 16274 22716
rect 16300 22439 16314 23257
rect 16294 22436 16320 22439
rect 16294 22407 16320 22410
rect 16340 21824 16366 21827
rect 16340 21795 16366 21798
rect 15834 21654 15860 21657
rect 15834 21625 15860 21628
rect 16156 21654 16182 21657
rect 16156 21625 16182 21628
rect 16248 21654 16274 21657
rect 16248 21625 16274 21628
rect 15840 20707 15854 21625
rect 16254 21385 16268 21625
rect 16248 21382 16274 21385
rect 16248 21353 16274 21356
rect 16248 21178 16274 21181
rect 16248 21149 16274 21152
rect 15794 20693 15854 20707
rect 15696 18934 15722 18937
rect 15696 18905 15722 18908
rect 15742 18934 15768 18937
rect 15742 18905 15768 18908
rect 15650 18900 15676 18903
rect 15650 18871 15676 18874
rect 15696 18832 15722 18835
rect 15696 18803 15722 18806
rect 15650 18662 15676 18665
rect 15650 18633 15676 18636
rect 15656 16965 15670 18633
rect 15702 18631 15716 18803
rect 15748 18733 15762 18905
rect 15742 18730 15768 18733
rect 15742 18701 15768 18704
rect 15794 18665 15808 20693
rect 15926 20464 15952 20467
rect 15926 20435 15952 20438
rect 15880 20294 15906 20297
rect 15880 20265 15906 20268
rect 15834 20226 15860 20229
rect 15834 20197 15860 20200
rect 15788 18662 15814 18665
rect 15788 18633 15814 18636
rect 15696 18628 15722 18631
rect 15696 18599 15722 18602
rect 15840 18563 15854 20197
rect 15886 19923 15900 20265
rect 15932 20195 15946 20435
rect 15926 20192 15952 20195
rect 15926 20163 15952 20166
rect 15972 20192 15998 20195
rect 15972 20163 15998 20166
rect 15880 19920 15906 19923
rect 15880 19891 15906 19894
rect 15742 18560 15768 18563
rect 15742 18531 15768 18534
rect 15788 18560 15814 18563
rect 15788 18531 15814 18534
rect 15834 18560 15860 18563
rect 15834 18531 15860 18534
rect 15748 18393 15762 18531
rect 15794 18461 15808 18531
rect 15788 18458 15814 18461
rect 15788 18429 15814 18432
rect 15742 18390 15768 18393
rect 15742 18361 15768 18364
rect 15650 16962 15676 16965
rect 15650 16933 15676 16936
rect 15834 16962 15860 16965
rect 15860 16942 15900 16956
rect 15834 16933 15860 16936
rect 15604 15160 15630 15163
rect 15604 15131 15630 15134
rect 15512 15126 15538 15129
rect 15472 15106 15512 15120
rect 15420 14616 15446 14619
rect 15420 14587 15446 14590
rect 15426 14117 15440 14587
rect 15472 14585 15486 15106
rect 15512 15097 15538 15100
rect 15466 14582 15492 14585
rect 15466 14553 15492 14556
rect 15656 14347 15670 16933
rect 15886 16769 15900 16942
rect 15932 16905 15946 20163
rect 15978 20025 15992 20163
rect 15972 20022 15998 20025
rect 15972 19993 15998 19996
rect 16110 20022 16136 20025
rect 16110 19993 16136 19996
rect 15972 19920 15998 19923
rect 15972 19891 15998 19894
rect 15978 19719 15992 19891
rect 16116 19719 16130 19993
rect 15972 19716 15998 19719
rect 15972 19687 15998 19690
rect 16110 19716 16136 19719
rect 16110 19687 16136 19690
rect 15978 18631 15992 19687
rect 16254 19685 16268 21149
rect 16346 21045 16360 21795
rect 16392 21181 16406 23971
rect 16714 23527 16728 24039
rect 17030 24000 17056 24003
rect 17030 23971 17056 23974
rect 16708 23524 16734 23527
rect 16708 23495 16734 23498
rect 16524 23286 16550 23289
rect 16524 23257 16550 23260
rect 16530 23085 16544 23257
rect 16570 23252 16596 23255
rect 16570 23223 16596 23226
rect 16524 23082 16550 23085
rect 16524 23053 16550 23056
rect 16530 22983 16544 23053
rect 16524 22980 16550 22983
rect 16524 22951 16550 22954
rect 16432 22946 16458 22949
rect 16432 22917 16458 22920
rect 16438 22507 16452 22917
rect 16432 22504 16458 22507
rect 16432 22475 16458 22478
rect 16438 22167 16452 22475
rect 16432 22164 16458 22167
rect 16432 22135 16458 22138
rect 16431 21944 16459 21948
rect 16431 21911 16459 21916
rect 16438 21827 16452 21911
rect 16432 21824 16458 21827
rect 16432 21795 16458 21798
rect 16524 21824 16550 21827
rect 16524 21795 16550 21798
rect 16432 21620 16458 21623
rect 16432 21591 16458 21594
rect 16386 21178 16412 21181
rect 16386 21149 16412 21152
rect 16340 21042 16366 21045
rect 16340 21013 16366 21016
rect 16248 19682 16274 19685
rect 16248 19653 16274 19656
rect 15972 18628 15998 18631
rect 15972 18599 15998 18602
rect 16156 18628 16182 18631
rect 16156 18599 16182 18602
rect 16202 18628 16228 18631
rect 16202 18599 16228 18602
rect 16162 18087 16176 18599
rect 16156 18084 16182 18087
rect 16156 18055 16182 18058
rect 16208 17475 16222 18599
rect 16202 17472 16228 17475
rect 16202 17443 16228 17446
rect 16017 16980 16045 16984
rect 16017 16947 16018 16952
rect 16044 16947 16045 16952
rect 16018 16933 16044 16936
rect 15932 16891 16038 16905
rect 15971 16776 15999 16780
rect 15840 16761 15946 16769
rect 15834 16758 15946 16761
rect 15860 16755 15946 16758
rect 15834 16729 15860 16732
rect 15880 16656 15906 16659
rect 15880 16627 15906 16630
rect 15788 15330 15814 15333
rect 15788 15301 15814 15304
rect 15794 14925 15808 15301
rect 15788 14922 15814 14925
rect 15788 14893 15814 14896
rect 15886 14823 15900 16627
rect 15932 16421 15946 16755
rect 15971 16743 15972 16748
rect 15998 16743 15999 16748
rect 15972 16729 15998 16732
rect 15926 16418 15952 16421
rect 15926 16389 15952 16392
rect 16024 15877 16038 16891
rect 16208 16455 16222 17443
rect 16202 16452 16228 16455
rect 16202 16423 16228 16426
rect 15978 15863 16038 15877
rect 15926 15466 15952 15469
rect 15926 15437 15952 15440
rect 15880 14820 15906 14823
rect 15880 14791 15906 14794
rect 15932 14729 15946 15437
rect 15978 15367 15992 15863
rect 16202 15670 16228 15673
rect 16254 15664 16268 19653
rect 16228 15650 16268 15664
rect 16202 15641 16228 15644
rect 16248 15568 16274 15571
rect 16248 15539 16274 15542
rect 16064 15398 16090 15401
rect 16064 15369 16090 15372
rect 16156 15398 16182 15401
rect 16156 15369 16182 15372
rect 15972 15364 15998 15367
rect 15972 15335 15998 15338
rect 15886 14715 15946 14729
rect 15650 14344 15676 14347
rect 15650 14315 15676 14318
rect 15426 14103 15486 14117
rect 15420 14038 15446 14041
rect 15420 14009 15446 14012
rect 15426 13837 15440 14009
rect 15420 13834 15446 13837
rect 15420 13805 15446 13808
rect 15373 13580 15401 13584
rect 15328 13562 15354 13565
rect 15373 13547 15401 13552
rect 15328 13533 15354 13536
rect 15281 12356 15309 12360
rect 15281 12323 15309 12328
rect 15472 11952 15486 14103
rect 15656 14041 15670 14315
rect 15650 14038 15676 14041
rect 15650 14009 15676 14012
rect 15604 13460 15630 13463
rect 15604 13431 15630 13434
rect 15610 12409 15624 13431
rect 15886 13293 15900 14715
rect 15926 13732 15952 13735
rect 15926 13703 15952 13706
rect 15880 13290 15906 13293
rect 15880 13261 15906 13264
rect 15696 12644 15722 12647
rect 15696 12615 15722 12618
rect 15604 12406 15630 12409
rect 15604 12377 15630 12380
rect 15702 12205 15716 12615
rect 15742 12576 15768 12579
rect 15742 12547 15768 12550
rect 15748 12443 15762 12547
rect 15742 12440 15768 12443
rect 15742 12411 15768 12414
rect 15696 12202 15722 12205
rect 15696 12173 15722 12176
rect 15932 12103 15946 13703
rect 15926 12100 15952 12103
rect 15926 12071 15952 12074
rect 15788 12066 15814 12069
rect 15788 12037 15814 12040
rect 15465 11948 15493 11952
rect 15794 11933 15808 12037
rect 15465 11915 15493 11920
rect 15788 11930 15814 11933
rect 15788 11901 15814 11904
rect 15742 10842 15768 10845
rect 15742 10813 15768 10816
rect 14730 10774 14756 10777
rect 14730 10745 14756 10748
rect 15144 10774 15170 10777
rect 15144 10745 15170 10748
rect 14040 10740 14066 10743
rect 14040 10711 14066 10714
rect 13948 10570 13974 10573
rect 13948 10541 13974 10544
rect 13672 10502 13698 10505
rect 13672 10473 13698 10476
rect 13856 10502 13882 10505
rect 13856 10473 13882 10476
rect 13948 10502 13974 10505
rect 13948 10473 13974 10476
rect 12384 10468 12410 10471
rect 12384 10439 12410 10442
rect 13902 10434 13928 10437
rect 13902 10405 13928 10408
rect 13908 9893 13922 10405
rect 13902 9890 13928 9893
rect 13902 9861 13928 9864
rect 13810 9176 13836 9179
rect 13810 9147 13836 9150
rect 13626 8802 13652 8805
rect 13626 8773 13652 8776
rect 13632 6663 13646 8773
rect 13718 7952 13744 7955
rect 13718 7923 13744 7926
rect 13724 7751 13738 7923
rect 13718 7748 13744 7751
rect 13718 7719 13744 7722
rect 13816 7003 13830 9147
rect 13856 8802 13882 8805
rect 13856 8773 13882 8776
rect 13862 8023 13876 8773
rect 13856 8020 13882 8023
rect 13856 7991 13882 7994
rect 13862 7751 13876 7991
rect 13856 7748 13882 7751
rect 13856 7719 13882 7722
rect 13810 7000 13836 7003
rect 13810 6971 13836 6974
rect 13764 6864 13790 6867
rect 13764 6835 13790 6838
rect 13770 6663 13784 6835
rect 13626 6660 13652 6663
rect 13626 6631 13652 6634
rect 13764 6660 13790 6663
rect 13764 6631 13790 6634
rect 13632 5337 13646 6631
rect 13626 5334 13652 5337
rect 13626 5305 13652 5308
rect 13954 3457 13968 10473
rect 14046 10403 14060 10711
rect 14776 10536 14802 10539
rect 14776 10507 14802 10510
rect 14408 10468 14434 10471
rect 14408 10439 14434 10442
rect 14316 10434 14342 10437
rect 14316 10405 14342 10408
rect 14040 10400 14066 10403
rect 14040 10371 14066 10374
rect 14046 10199 14060 10371
rect 14322 10301 14336 10405
rect 14316 10298 14342 10301
rect 14316 10269 14342 10272
rect 14040 10196 14066 10199
rect 14040 10167 14066 10170
rect 14046 9383 14060 10167
rect 14414 9927 14428 10439
rect 14592 10434 14618 10437
rect 14592 10405 14618 10408
rect 14408 9924 14434 9927
rect 14408 9895 14434 9898
rect 14414 9757 14428 9895
rect 14598 9893 14612 10405
rect 14782 10267 14796 10507
rect 14868 10400 14894 10403
rect 14868 10371 14894 10374
rect 14776 10264 14802 10267
rect 14776 10235 14802 10238
rect 14874 10131 14888 10371
rect 14638 10128 14664 10131
rect 14638 10099 14664 10102
rect 14868 10128 14894 10131
rect 14868 10099 14894 10102
rect 14644 9927 14658 10099
rect 15098 9958 15124 9961
rect 15098 9929 15124 9932
rect 14638 9924 14664 9927
rect 14638 9895 14664 9898
rect 14592 9890 14618 9893
rect 14592 9861 14618 9864
rect 14408 9754 14434 9757
rect 14408 9725 14434 9728
rect 14362 9584 14388 9587
rect 14362 9555 14388 9558
rect 14368 9383 14382 9555
rect 14414 9383 14428 9725
rect 14500 9686 14526 9689
rect 14500 9657 14526 9660
rect 14040 9380 14066 9383
rect 14040 9351 14066 9354
rect 14362 9380 14388 9383
rect 14362 9351 14388 9354
rect 14408 9380 14434 9383
rect 14408 9351 14434 9354
rect 14046 8771 14060 9351
rect 14414 9179 14428 9351
rect 14506 9213 14520 9657
rect 14546 9312 14572 9315
rect 14546 9283 14572 9286
rect 14500 9210 14526 9213
rect 14500 9181 14526 9184
rect 14408 9176 14434 9179
rect 14408 9147 14434 9150
rect 14132 9142 14158 9145
rect 14132 9113 14158 9116
rect 14138 8907 14152 9113
rect 14414 8949 14428 9147
rect 14552 9145 14566 9283
rect 14644 9179 14658 9895
rect 15052 9720 15078 9723
rect 15052 9691 15078 9694
rect 15058 9485 15072 9691
rect 15052 9482 15078 9485
rect 15052 9453 15078 9456
rect 15104 9417 15118 9929
rect 15236 9856 15262 9859
rect 15236 9827 15262 9830
rect 15098 9414 15124 9417
rect 15098 9385 15124 9388
rect 14638 9176 14664 9179
rect 14638 9147 14664 9150
rect 14546 9142 14572 9145
rect 14506 9122 14546 9136
rect 14454 9040 14480 9043
rect 14454 9011 14480 9014
rect 14322 8935 14428 8949
rect 14460 8941 14474 9011
rect 14454 8938 14480 8941
rect 14132 8904 14158 8907
rect 14132 8875 14158 8878
rect 14322 8839 14336 8935
rect 14454 8909 14480 8912
rect 14408 8904 14434 8907
rect 14408 8875 14434 8878
rect 14316 8836 14342 8839
rect 14316 8807 14342 8810
rect 14040 8768 14066 8771
rect 14040 8739 14066 8742
rect 14414 8057 14428 8875
rect 14506 8057 14520 9122
rect 14546 9113 14572 9116
rect 14546 9074 14572 9077
rect 14546 9045 14572 9048
rect 14552 8057 14566 9045
rect 15104 8839 15118 9385
rect 15098 8836 15124 8839
rect 15098 8807 15124 8810
rect 15242 8805 15256 9827
rect 15466 9346 15492 9349
rect 15466 9317 15492 9320
rect 15472 9111 15486 9317
rect 15466 9108 15492 9111
rect 15466 9079 15492 9082
rect 15236 8802 15262 8805
rect 15236 8773 15262 8776
rect 15696 8802 15722 8805
rect 15696 8773 15722 8776
rect 14408 8054 14434 8057
rect 14408 8025 14434 8028
rect 14500 8054 14526 8057
rect 14500 8025 14526 8028
rect 14546 8054 14572 8057
rect 14546 8025 14572 8028
rect 14040 7782 14066 7785
rect 14040 7753 14066 7756
rect 14046 7241 14060 7753
rect 14414 7717 14428 8025
rect 14506 7819 14520 8025
rect 14500 7816 14526 7819
rect 14500 7787 14526 7790
rect 14552 7751 14566 8025
rect 14546 7748 14572 7751
rect 14546 7719 14572 7722
rect 14408 7714 14434 7717
rect 14408 7685 14434 7688
rect 14316 7476 14342 7479
rect 14316 7447 14342 7450
rect 14322 7309 14336 7447
rect 14316 7306 14342 7309
rect 14316 7277 14342 7280
rect 14040 7238 14066 7241
rect 14040 7209 14066 7212
rect 14322 7045 14336 7277
rect 14408 7204 14434 7207
rect 14408 7175 14434 7178
rect 14276 7031 14336 7045
rect 14276 6969 14290 7031
rect 14270 6966 14296 6969
rect 14270 6937 14296 6940
rect 14414 6901 14428 7175
rect 14408 6898 14434 6901
rect 14408 6869 14434 6872
rect 14414 6765 14428 6869
rect 14408 6762 14434 6765
rect 14408 6733 14434 6736
rect 15242 5541 15256 8773
rect 15702 8125 15716 8773
rect 15696 8122 15722 8125
rect 15696 8093 15722 8096
rect 15748 8065 15762 10813
rect 15794 10471 15808 11901
rect 15978 11865 15992 15335
rect 16018 15024 16044 15027
rect 16018 14995 16044 14998
rect 16024 14857 16038 14995
rect 16018 14854 16044 14857
rect 16018 14825 16044 14828
rect 16070 14755 16084 15369
rect 16110 15364 16136 15367
rect 16110 15335 16136 15338
rect 16064 14752 16090 14755
rect 16064 14723 16090 14726
rect 16018 13494 16044 13497
rect 16018 13465 16044 13468
rect 16024 13293 16038 13465
rect 16018 13290 16044 13293
rect 16018 13261 16044 13264
rect 16116 12171 16130 15335
rect 16162 14789 16176 15369
rect 16254 15333 16268 15539
rect 16346 15333 16360 21013
rect 16438 15469 16452 21591
rect 16530 18393 16544 21795
rect 16576 21113 16590 23223
rect 16714 22983 16728 23495
rect 16708 22980 16734 22983
rect 16708 22951 16734 22954
rect 16616 22436 16642 22439
rect 16616 22407 16642 22410
rect 16622 22235 16636 22407
rect 16616 22232 16642 22235
rect 16616 22203 16642 22206
rect 16622 21895 16636 22203
rect 16714 22099 16728 22951
rect 16708 22096 16734 22099
rect 16708 22067 16734 22070
rect 16616 21892 16642 21895
rect 16616 21863 16642 21866
rect 16622 21453 16636 21863
rect 16714 21691 16728 22067
rect 16708 21688 16734 21691
rect 16708 21659 16734 21662
rect 16616 21450 16642 21453
rect 16616 21421 16642 21424
rect 16714 21351 16728 21659
rect 16708 21348 16734 21351
rect 16708 21319 16734 21322
rect 16570 21110 16596 21113
rect 16570 21081 16596 21084
rect 17036 20467 17050 23971
rect 17082 23561 17096 24583
rect 17128 24105 17142 24787
rect 17266 24649 17280 24889
rect 17260 24646 17286 24649
rect 17260 24617 17286 24620
rect 17122 24102 17148 24105
rect 17122 24073 17148 24076
rect 17076 23558 17102 23561
rect 17076 23529 17102 23532
rect 17082 23433 17096 23529
rect 17266 23493 17280 24617
rect 17260 23490 17286 23493
rect 17260 23461 17286 23464
rect 17082 23419 17188 23433
rect 17122 23354 17148 23357
rect 17122 23325 17148 23328
rect 17128 22832 17142 23325
rect 17174 23289 17188 23419
rect 17266 23323 17280 23461
rect 17260 23320 17286 23323
rect 17260 23291 17286 23294
rect 17168 23286 17194 23289
rect 17168 23257 17194 23260
rect 17121 22828 17149 22832
rect 17121 22795 17149 22800
rect 17030 20464 17056 20467
rect 17030 20435 17056 20438
rect 16892 20294 16918 20297
rect 16892 20265 16918 20268
rect 16524 18390 16550 18393
rect 16524 18361 16550 18364
rect 16478 18050 16504 18053
rect 16478 18021 16504 18024
rect 16484 16984 16498 18021
rect 16477 16980 16505 16984
rect 16477 16947 16505 16952
rect 16530 16693 16544 18361
rect 16524 16690 16550 16693
rect 16524 16661 16550 16664
rect 16432 15466 16458 15469
rect 16432 15437 16458 15440
rect 16898 15367 16912 20265
rect 17036 20186 17050 20435
rect 17076 20192 17102 20195
rect 17036 20172 17076 20186
rect 17076 20163 17102 20166
rect 17128 18393 17142 22795
rect 17174 22235 17188 23257
rect 17398 22946 17424 22949
rect 17398 22917 17424 22920
rect 17168 22232 17194 22235
rect 17168 22203 17194 22206
rect 17404 22133 17418 22917
rect 17398 22130 17424 22133
rect 17398 22101 17424 22104
rect 17404 21657 17418 22101
rect 17398 21654 17424 21657
rect 17398 21625 17424 21628
rect 17404 21351 17418 21625
rect 17398 21348 17424 21351
rect 17398 21319 17424 21322
rect 17260 21144 17286 21147
rect 17260 21115 17286 21118
rect 17214 21110 17240 21113
rect 17214 21081 17240 21084
rect 17168 21042 17194 21045
rect 17168 21013 17194 21016
rect 17174 20297 17188 21013
rect 17168 20294 17194 20297
rect 17168 20265 17194 20268
rect 17220 20263 17234 21081
rect 17214 20260 17240 20263
rect 17214 20231 17240 20234
rect 17168 18560 17194 18563
rect 17168 18531 17194 18534
rect 17174 18461 17188 18531
rect 17168 18458 17194 18461
rect 17168 18429 17194 18432
rect 17266 18393 17280 21115
rect 17306 20260 17332 20263
rect 17306 20231 17332 20234
rect 17398 20260 17424 20263
rect 17398 20231 17424 20234
rect 17312 20025 17326 20231
rect 17306 20022 17332 20025
rect 17306 19993 17332 19996
rect 17404 19821 17418 20231
rect 17398 19818 17424 19821
rect 17398 19789 17424 19792
rect 17122 18390 17148 18393
rect 17122 18361 17148 18364
rect 17214 18390 17240 18393
rect 17214 18361 17240 18364
rect 17260 18390 17286 18393
rect 17260 18361 17286 18364
rect 17030 17268 17056 17271
rect 17030 17239 17056 17242
rect 16938 15466 16964 15469
rect 16938 15437 16964 15440
rect 16944 15367 16958 15437
rect 16892 15364 16918 15367
rect 16892 15335 16918 15338
rect 16938 15364 16964 15367
rect 16938 15335 16964 15338
rect 16202 15330 16228 15333
rect 16202 15301 16228 15304
rect 16248 15330 16274 15333
rect 16248 15301 16274 15304
rect 16340 15330 16366 15333
rect 16340 15301 16366 15304
rect 16386 15330 16412 15333
rect 16386 15301 16412 15304
rect 16570 15330 16596 15333
rect 16570 15301 16596 15304
rect 16156 14786 16182 14789
rect 16156 14757 16182 14760
rect 16208 14483 16222 15301
rect 16202 14480 16228 14483
rect 16202 14451 16228 14454
rect 16293 13648 16321 13652
rect 16293 13615 16321 13620
rect 16300 13565 16314 13615
rect 16294 13562 16320 13565
rect 16294 13533 16320 13536
rect 16300 13191 16314 13533
rect 16294 13188 16320 13191
rect 16294 13159 16320 13162
rect 16294 12610 16320 12613
rect 16294 12581 16320 12584
rect 16300 12307 16314 12581
rect 16346 12477 16360 15301
rect 16392 15197 16406 15301
rect 16386 15194 16412 15197
rect 16386 15165 16412 15168
rect 16576 14925 16590 15301
rect 16570 14922 16596 14925
rect 16570 14893 16596 14896
rect 16754 14038 16780 14041
rect 16754 14009 16780 14012
rect 16760 13837 16774 14009
rect 16944 14007 16958 15335
rect 17036 15324 17050 17239
rect 17128 16999 17142 18361
rect 17220 18189 17234 18361
rect 17214 18186 17240 18189
rect 17214 18157 17240 18160
rect 17122 16996 17148 16999
rect 17122 16967 17148 16970
rect 17168 16996 17194 16999
rect 17168 16967 17194 16970
rect 17076 16928 17102 16931
rect 17076 16899 17102 16902
rect 17082 16795 17096 16899
rect 17076 16792 17102 16795
rect 17076 16763 17102 16766
rect 17122 16758 17148 16761
rect 17122 16729 17148 16732
rect 17128 16712 17142 16729
rect 17121 16708 17149 16712
rect 17121 16675 17149 16680
rect 17174 16557 17188 16967
rect 17266 16795 17280 18361
rect 17306 16928 17332 16931
rect 17306 16899 17332 16902
rect 17260 16792 17286 16795
rect 17260 16763 17286 16766
rect 17214 16656 17240 16659
rect 17214 16627 17240 16630
rect 17168 16554 17194 16557
rect 17168 16525 17194 16528
rect 17220 16455 17234 16627
rect 17312 16455 17326 16899
rect 17214 16452 17240 16455
rect 17214 16423 17240 16426
rect 17306 16452 17332 16455
rect 17306 16423 17332 16426
rect 17260 16384 17286 16387
rect 17260 16355 17286 16358
rect 17168 15330 17194 15333
rect 17036 15310 17168 15324
rect 17168 15301 17194 15304
rect 17174 14381 17188 15301
rect 17168 14378 17194 14381
rect 17168 14349 17194 14352
rect 17214 14208 17240 14211
rect 17214 14179 17240 14182
rect 16938 14004 16964 14007
rect 16938 13975 16964 13978
rect 17076 14004 17102 14007
rect 17076 13975 17102 13978
rect 16754 13834 16780 13837
rect 16754 13805 16780 13808
rect 17082 13769 17096 13975
rect 16800 13766 16826 13769
rect 16800 13737 16826 13740
rect 17076 13766 17102 13769
rect 17076 13737 17102 13740
rect 16524 13392 16550 13395
rect 16524 13363 16550 13366
rect 16432 12984 16458 12987
rect 16432 12955 16458 12958
rect 16438 12647 16452 12955
rect 16478 12950 16504 12953
rect 16478 12921 16504 12924
rect 16432 12644 16458 12647
rect 16432 12615 16458 12618
rect 16484 12613 16498 12921
rect 16530 12647 16544 13363
rect 16570 13188 16596 13191
rect 16570 13159 16596 13162
rect 16576 12919 16590 13159
rect 16570 12916 16596 12919
rect 16570 12887 16596 12890
rect 16570 12678 16596 12681
rect 16570 12649 16596 12652
rect 16524 12644 16550 12647
rect 16524 12615 16550 12618
rect 16478 12610 16504 12613
rect 16478 12581 16504 12584
rect 16340 12474 16366 12477
rect 16340 12445 16366 12448
rect 16294 12304 16320 12307
rect 16294 12275 16320 12278
rect 16110 12168 16136 12171
rect 16110 12139 16136 12142
rect 16110 12100 16136 12103
rect 16110 12071 16136 12074
rect 15972 11862 15998 11865
rect 15972 11833 15998 11836
rect 16116 11491 16130 12071
rect 16300 12069 16314 12275
rect 16294 12066 16320 12069
rect 16294 12037 16320 12040
rect 16386 11896 16412 11899
rect 16386 11867 16412 11870
rect 16248 11862 16274 11865
rect 16248 11833 16274 11836
rect 16340 11862 16366 11865
rect 16340 11833 16366 11836
rect 16110 11488 16136 11491
rect 16110 11459 16136 11462
rect 16254 11465 16268 11833
rect 16346 11559 16360 11833
rect 16392 11559 16406 11867
rect 16530 11865 16544 12615
rect 16576 12069 16590 12649
rect 16806 12205 16820 13737
rect 17082 13531 17096 13737
rect 17076 13528 17102 13531
rect 17076 13499 17102 13502
rect 16938 13222 16964 13225
rect 16938 13193 16964 13196
rect 16800 12202 16826 12205
rect 16800 12173 16826 12176
rect 16570 12066 16596 12069
rect 16570 12037 16596 12040
rect 16524 11862 16550 11865
rect 16524 11833 16550 11836
rect 16340 11556 16366 11559
rect 16340 11527 16366 11530
rect 16386 11556 16412 11559
rect 16386 11527 16412 11530
rect 15880 10944 15906 10947
rect 15880 10915 15906 10918
rect 15788 10468 15814 10471
rect 15788 10439 15814 10442
rect 15886 10267 15900 10915
rect 15972 10434 15998 10437
rect 15972 10405 15998 10408
rect 15880 10264 15906 10267
rect 15880 10235 15906 10238
rect 15978 10199 15992 10405
rect 15972 10196 15998 10199
rect 15972 10167 15998 10170
rect 15978 9995 15992 10167
rect 15972 9992 15998 9995
rect 15972 9963 15998 9966
rect 15788 9312 15814 9315
rect 15880 9312 15906 9315
rect 15814 9292 15854 9306
rect 15788 9283 15814 9286
rect 15840 8839 15854 9292
rect 15880 9283 15906 9286
rect 15788 8836 15814 8839
rect 15788 8807 15814 8810
rect 15834 8836 15860 8839
rect 15834 8807 15860 8810
rect 15702 8051 15762 8065
rect 15702 6217 15716 8051
rect 15794 7581 15808 8807
rect 15886 8023 15900 9283
rect 15978 9221 15992 9963
rect 16116 9383 16130 11459
rect 16254 11451 16360 11465
rect 16156 11318 16182 11321
rect 16156 11289 16182 11292
rect 16162 11015 16176 11289
rect 16248 11250 16274 11253
rect 16248 11221 16274 11224
rect 16202 11216 16228 11219
rect 16202 11187 16228 11190
rect 16156 11012 16182 11015
rect 16156 10983 16182 10986
rect 16208 10505 16222 11187
rect 16254 11015 16268 11221
rect 16346 11219 16360 11451
rect 16340 11216 16366 11219
rect 16340 11187 16366 11190
rect 16346 11049 16360 11187
rect 16340 11046 16366 11049
rect 16340 11017 16366 11020
rect 16392 11015 16406 11527
rect 16576 11321 16590 12037
rect 16662 12032 16688 12035
rect 16662 12003 16688 12006
rect 16668 11593 16682 12003
rect 16662 11590 16688 11593
rect 16662 11561 16688 11564
rect 16570 11318 16596 11321
rect 16570 11289 16596 11292
rect 16248 11012 16274 11015
rect 16248 10983 16274 10986
rect 16386 11012 16412 11015
rect 16386 10983 16412 10986
rect 16524 10842 16550 10845
rect 16524 10813 16550 10816
rect 16202 10502 16228 10505
rect 16202 10473 16228 10476
rect 16530 10437 16544 10813
rect 16248 10434 16274 10437
rect 16248 10405 16274 10408
rect 16524 10434 16550 10437
rect 16524 10405 16550 10408
rect 16254 10267 16268 10405
rect 16248 10264 16274 10267
rect 16248 10235 16274 10238
rect 16944 9655 16958 13193
rect 17168 13120 17194 13123
rect 17168 13091 17194 13094
rect 17076 12916 17102 12919
rect 17076 12887 17102 12890
rect 17082 12443 17096 12887
rect 17174 12579 17188 13091
rect 17168 12576 17194 12579
rect 17168 12547 17194 12550
rect 17076 12440 17102 12443
rect 17076 12411 17102 12414
rect 17174 12409 17188 12547
rect 17220 12417 17234 14179
rect 17266 14075 17280 16355
rect 17260 14072 17286 14075
rect 17260 14043 17286 14046
rect 17450 12987 17464 27779
rect 17680 27675 17694 27847
rect 17910 27811 17924 28119
rect 18094 28117 18108 28153
rect 18088 28114 18114 28117
rect 18088 28085 18114 28088
rect 18094 27879 18108 28085
rect 18088 27876 18114 27879
rect 18088 27847 18114 27850
rect 17904 27808 17930 27811
rect 17904 27779 17930 27782
rect 17674 27672 17700 27675
rect 17674 27643 17700 27646
rect 17996 27638 18022 27641
rect 17996 27609 18022 27612
rect 18002 27165 18016 27609
rect 18094 27573 18108 27847
rect 18456 27638 18482 27641
rect 18456 27609 18482 27612
rect 18088 27570 18114 27573
rect 18088 27541 18114 27544
rect 18364 27570 18390 27573
rect 18364 27541 18390 27544
rect 17996 27162 18022 27165
rect 17996 27133 18022 27136
rect 18370 27063 18384 27541
rect 18226 27060 18252 27063
rect 18226 27031 18252 27034
rect 18272 27060 18298 27063
rect 18272 27031 18298 27034
rect 18364 27060 18390 27063
rect 18364 27031 18390 27034
rect 17812 26788 17838 26791
rect 17812 26759 17838 26762
rect 17674 26754 17700 26757
rect 17674 26725 17700 26728
rect 17490 26210 17516 26213
rect 17490 26181 17516 26184
rect 17496 25805 17510 26181
rect 17680 26179 17694 26725
rect 17766 26720 17792 26723
rect 17766 26691 17792 26694
rect 17720 26516 17746 26519
rect 17720 26487 17746 26490
rect 17726 26213 17740 26487
rect 17720 26210 17746 26213
rect 17720 26181 17746 26184
rect 17674 26176 17700 26179
rect 17674 26147 17700 26150
rect 17490 25802 17516 25805
rect 17490 25773 17516 25776
rect 17720 25122 17746 25125
rect 17720 25093 17746 25096
rect 17726 24377 17740 25093
rect 17772 24445 17786 26691
rect 17818 26621 17832 26759
rect 17904 26720 17930 26723
rect 17904 26691 17930 26694
rect 17812 26618 17838 26621
rect 17812 26589 17838 26592
rect 17910 26519 17924 26691
rect 18042 26550 18068 26553
rect 18002 26530 18042 26544
rect 17904 26516 17930 26519
rect 17904 26487 17930 26490
rect 17858 26448 17884 26451
rect 17858 26419 17884 26422
rect 17864 26349 17878 26419
rect 17858 26346 17884 26349
rect 17858 26317 17884 26320
rect 18002 26315 18016 26530
rect 18042 26521 18068 26524
rect 17996 26312 18022 26315
rect 17996 26283 18022 26286
rect 17950 26210 17976 26213
rect 17950 26181 17976 26184
rect 17956 26043 17970 26181
rect 18002 26179 18016 26283
rect 17996 26176 18022 26179
rect 17996 26147 18022 26150
rect 17950 26040 17976 26043
rect 17950 26011 17976 26014
rect 17904 25462 17930 25465
rect 17904 25433 17930 25436
rect 17910 24615 17924 25433
rect 17904 24612 17930 24615
rect 17904 24583 17930 24586
rect 17766 24442 17792 24445
rect 17766 24413 17792 24416
rect 17720 24374 17746 24377
rect 17720 24345 17746 24348
rect 17536 24340 17562 24343
rect 17536 24311 17562 24314
rect 17542 23085 17556 24311
rect 17910 24071 17924 24583
rect 17904 24068 17930 24071
rect 17904 24039 17930 24042
rect 17910 23901 17924 24039
rect 18002 24003 18016 26147
rect 18232 24717 18246 27031
rect 18278 26893 18292 27031
rect 18272 26890 18298 26893
rect 18272 26861 18298 26864
rect 18462 26825 18476 27609
rect 18456 26822 18482 26825
rect 18456 26793 18482 26796
rect 18508 26612 18522 28357
rect 19008 28182 19034 28185
rect 19008 28153 19034 28156
rect 18686 28148 18712 28151
rect 18686 28119 18712 28122
rect 18692 27879 18706 28119
rect 18686 27876 18712 27879
rect 18686 27847 18712 27850
rect 18732 27842 18758 27845
rect 18732 27813 18758 27816
rect 18738 27437 18752 27813
rect 19014 27811 19028 28153
rect 19244 28083 19258 28425
rect 19376 28420 19402 28423
rect 19376 28391 19402 28394
rect 19382 28253 19396 28391
rect 19376 28250 19402 28253
rect 19376 28221 19402 28224
rect 20164 28151 20178 28663
rect 20302 28525 20316 28663
rect 20296 28522 20322 28525
rect 20296 28493 20322 28496
rect 20158 28148 20184 28151
rect 20158 28119 20184 28122
rect 20342 28148 20368 28151
rect 20342 28119 20368 28122
rect 19238 28080 19264 28083
rect 19238 28051 19264 28054
rect 19100 27876 19126 27879
rect 19100 27847 19126 27850
rect 19008 27808 19034 27811
rect 19008 27779 19034 27782
rect 19014 27641 19028 27779
rect 19008 27638 19034 27641
rect 19008 27609 19034 27612
rect 18778 27570 18804 27573
rect 18778 27541 18804 27544
rect 18732 27434 18758 27437
rect 18732 27405 18758 27408
rect 18784 27369 18798 27541
rect 18778 27366 18804 27369
rect 18778 27337 18804 27340
rect 19106 27335 19120 27847
rect 19244 27675 19258 28051
rect 19468 27808 19494 27811
rect 19468 27779 19494 27782
rect 19238 27672 19264 27675
rect 19238 27643 19264 27646
rect 19376 27536 19402 27539
rect 19376 27507 19402 27510
rect 19100 27332 19126 27335
rect 19100 27303 19126 27306
rect 19106 26791 19120 27303
rect 19382 27301 19396 27507
rect 19474 27437 19488 27779
rect 19468 27434 19494 27437
rect 19468 27405 19494 27408
rect 19422 27332 19448 27335
rect 19422 27303 19448 27306
rect 19376 27298 19402 27301
rect 19376 27269 19402 27272
rect 19100 26788 19126 26791
rect 19100 26759 19126 26762
rect 18640 26754 18666 26757
rect 18640 26725 18666 26728
rect 18462 26598 18522 26612
rect 18318 25496 18344 25499
rect 18318 25467 18344 25470
rect 18324 24989 18338 25467
rect 18364 25190 18390 25193
rect 18364 25161 18390 25164
rect 18318 24986 18344 24989
rect 18318 24957 18344 24960
rect 18324 24887 18338 24957
rect 18318 24884 18344 24887
rect 18318 24855 18344 24858
rect 18226 24714 18252 24717
rect 18226 24685 18252 24688
rect 18088 24068 18114 24071
rect 18088 24039 18114 24042
rect 17996 24000 18022 24003
rect 17996 23971 18022 23974
rect 17904 23898 17930 23901
rect 17904 23869 17930 23872
rect 17910 23595 17924 23869
rect 18094 23799 18108 24039
rect 18370 23833 18384 25161
rect 18462 24887 18476 26598
rect 18502 26550 18528 26553
rect 18502 26521 18528 26524
rect 18508 26077 18522 26521
rect 18646 26436 18660 26725
rect 19106 26485 19120 26759
rect 19382 26757 19396 27269
rect 19376 26754 19402 26757
rect 19376 26725 19402 26728
rect 19100 26482 19126 26485
rect 19100 26453 19126 26456
rect 18639 26432 18667 26436
rect 18639 26399 18667 26404
rect 18870 26278 18896 26281
rect 18870 26249 18896 26252
rect 18640 26210 18666 26213
rect 18640 26181 18666 26184
rect 18502 26074 18528 26077
rect 18502 26045 18528 26048
rect 18502 25972 18528 25975
rect 18502 25943 18528 25946
rect 18508 25193 18522 25943
rect 18502 25190 18528 25193
rect 18502 25161 18528 25164
rect 18548 25122 18574 25125
rect 18548 25093 18574 25096
rect 18554 24921 18568 25093
rect 18548 24918 18574 24921
rect 18548 24889 18574 24892
rect 18456 24884 18482 24887
rect 18456 24855 18482 24858
rect 18462 24181 18476 24855
rect 18554 24615 18568 24889
rect 18594 24646 18620 24649
rect 18594 24617 18620 24620
rect 18548 24612 18574 24615
rect 18548 24583 18574 24586
rect 18462 24167 18568 24181
rect 18456 24136 18482 24139
rect 18456 24107 18482 24110
rect 18462 23867 18476 24107
rect 18502 24034 18528 24037
rect 18502 24005 18528 24008
rect 18456 23864 18482 23867
rect 18456 23835 18482 23838
rect 18364 23830 18390 23833
rect 18364 23801 18390 23804
rect 17950 23796 17976 23799
rect 17950 23767 17976 23770
rect 18088 23796 18114 23799
rect 18088 23767 18114 23770
rect 17904 23592 17930 23595
rect 17904 23563 17930 23566
rect 17812 23490 17838 23493
rect 17812 23461 17838 23464
rect 17536 23082 17562 23085
rect 17536 23053 17562 23056
rect 17674 23014 17700 23017
rect 17674 22985 17700 22988
rect 17490 22980 17516 22983
rect 17490 22951 17516 22954
rect 17582 22980 17608 22983
rect 17582 22951 17608 22954
rect 17496 22779 17510 22951
rect 17490 22776 17516 22779
rect 17490 22747 17516 22750
rect 17496 22439 17510 22747
rect 17490 22436 17516 22439
rect 17490 22407 17516 22410
rect 17496 21997 17510 22407
rect 17588 22371 17602 22951
rect 17628 22708 17654 22711
rect 17628 22679 17654 22682
rect 17634 22507 17648 22679
rect 17680 22634 17694 22985
rect 17818 22983 17832 23461
rect 17910 23289 17924 23563
rect 17956 23561 17970 23767
rect 17950 23558 17976 23561
rect 17950 23529 17976 23532
rect 18134 23558 18160 23561
rect 18134 23529 18160 23532
rect 17950 23456 17976 23459
rect 17950 23427 17976 23430
rect 17956 23357 17970 23427
rect 17950 23354 17976 23357
rect 17950 23325 17976 23328
rect 18140 23289 18154 23529
rect 17904 23286 17930 23289
rect 17904 23257 17930 23260
rect 18134 23286 18160 23289
rect 18134 23257 18160 23260
rect 17812 22980 17838 22983
rect 17812 22951 17838 22954
rect 17818 22779 17832 22951
rect 17910 22949 17924 23257
rect 17904 22946 17930 22949
rect 17904 22917 17930 22920
rect 17950 22912 17976 22915
rect 17950 22883 17976 22886
rect 17812 22776 17838 22779
rect 17812 22747 17838 22750
rect 17766 22742 17792 22745
rect 17766 22713 17792 22716
rect 17720 22640 17746 22643
rect 17680 22620 17720 22634
rect 17628 22504 17654 22507
rect 17628 22475 17654 22478
rect 17680 22473 17694 22620
rect 17720 22611 17746 22614
rect 17772 22541 17786 22713
rect 17766 22538 17792 22541
rect 17766 22509 17792 22512
rect 17674 22470 17700 22473
rect 17674 22441 17700 22444
rect 17582 22368 17608 22371
rect 17582 22339 17608 22342
rect 17536 22232 17562 22235
rect 17536 22203 17562 22206
rect 17490 21994 17516 21997
rect 17490 21965 17516 21968
rect 17542 21895 17556 22203
rect 17536 21892 17562 21895
rect 17536 21863 17562 21866
rect 17680 17271 17694 22441
rect 17766 22368 17792 22371
rect 17766 22339 17792 22342
rect 17772 22167 17786 22339
rect 17818 22201 17832 22747
rect 17904 22742 17930 22745
rect 17904 22713 17930 22716
rect 17910 22541 17924 22713
rect 17904 22538 17930 22541
rect 17904 22509 17930 22512
rect 17910 22235 17924 22509
rect 17956 22439 17970 22883
rect 18370 22473 18384 23801
rect 18508 23629 18522 24005
rect 18502 23626 18528 23629
rect 18502 23597 18528 23600
rect 18554 23561 18568 24167
rect 18600 24071 18614 24617
rect 18646 24105 18660 26181
rect 18876 25533 18890 26249
rect 19106 26247 19120 26453
rect 19382 26247 19396 26725
rect 19100 26244 19126 26247
rect 19100 26215 19126 26218
rect 19376 26244 19402 26247
rect 19376 26215 19402 26218
rect 19106 25975 19120 26215
rect 19100 25972 19126 25975
rect 19100 25943 19126 25946
rect 19428 25537 19442 27303
rect 20164 27063 20178 28119
rect 20348 27981 20362 28119
rect 20342 27978 20368 27981
rect 20342 27949 20368 27952
rect 20158 27060 20184 27063
rect 20158 27031 20184 27034
rect 20296 27060 20322 27063
rect 20296 27031 20322 27034
rect 20434 27060 20460 27063
rect 20434 27031 20460 27034
rect 20250 26550 20276 26553
rect 20250 26521 20276 26524
rect 20256 26043 20270 26521
rect 20302 26485 20316 27031
rect 20440 26621 20454 27031
rect 20434 26618 20460 26621
rect 20434 26589 20460 26592
rect 20296 26482 20322 26485
rect 20296 26453 20322 26456
rect 20250 26040 20276 26043
rect 20250 26011 20276 26014
rect 18870 25530 18896 25533
rect 19428 25523 19488 25537
rect 18870 25501 18896 25504
rect 18778 25462 18804 25465
rect 18778 25433 18804 25436
rect 18686 25088 18712 25091
rect 18686 25059 18712 25062
rect 18692 24887 18706 25059
rect 18686 24884 18712 24887
rect 18686 24855 18712 24858
rect 18784 24853 18798 25433
rect 18916 25428 18942 25431
rect 18916 25399 18942 25402
rect 18922 24887 18936 25399
rect 19100 25360 19126 25363
rect 19100 25331 19126 25334
rect 19106 25159 19120 25331
rect 19100 25156 19126 25159
rect 19100 25127 19126 25130
rect 18916 24884 18942 24887
rect 18916 24855 18942 24858
rect 18778 24850 18804 24853
rect 18778 24821 18804 24824
rect 19422 24646 19448 24649
rect 19422 24617 19448 24620
rect 18640 24102 18666 24105
rect 18640 24073 18666 24076
rect 18594 24068 18620 24071
rect 18594 24039 18620 24042
rect 18594 24000 18620 24003
rect 18594 23971 18620 23974
rect 18548 23558 18574 23561
rect 18548 23529 18574 23532
rect 18502 23286 18528 23289
rect 18502 23257 18528 23260
rect 18508 23051 18522 23257
rect 18410 23048 18436 23051
rect 18410 23019 18436 23022
rect 18502 23048 18528 23051
rect 18502 23019 18528 23022
rect 18364 22470 18390 22473
rect 18364 22441 18390 22444
rect 17950 22436 17976 22439
rect 17950 22407 17976 22410
rect 17904 22232 17930 22235
rect 17904 22203 17930 22206
rect 17812 22198 17838 22201
rect 17812 22169 17838 22172
rect 17766 22164 17792 22167
rect 17766 22135 17792 22138
rect 17720 21926 17746 21929
rect 17720 21897 17746 21900
rect 17726 21691 17740 21897
rect 17818 21895 17832 22169
rect 17904 21926 17930 21929
rect 17904 21897 17930 21900
rect 17812 21892 17838 21895
rect 17812 21863 17838 21866
rect 17720 21688 17746 21691
rect 17720 21659 17746 21662
rect 17910 21623 17924 21897
rect 18226 21722 18252 21725
rect 18226 21693 18252 21696
rect 17904 21620 17930 21623
rect 17904 21591 17930 21594
rect 18232 21147 18246 21693
rect 18226 21144 18252 21147
rect 18226 21115 18252 21118
rect 17996 20906 18022 20909
rect 17996 20877 18022 20880
rect 17858 20022 17884 20025
rect 17858 19993 17884 19996
rect 17720 19988 17746 19991
rect 17720 19959 17746 19962
rect 17726 19277 17740 19959
rect 17864 19285 17878 19993
rect 17720 19274 17746 19277
rect 17864 19271 17970 19285
rect 17720 19245 17746 19248
rect 17726 18937 17740 19245
rect 17956 19107 17970 19271
rect 17950 19104 17976 19107
rect 17950 19075 17976 19078
rect 17956 18937 17970 19075
rect 17720 18934 17746 18937
rect 17720 18905 17746 18908
rect 17950 18934 17976 18937
rect 17950 18905 17976 18908
rect 17726 18087 17740 18905
rect 17956 18393 17970 18905
rect 17950 18390 17976 18393
rect 17950 18361 17976 18364
rect 17720 18084 17746 18087
rect 17720 18055 17746 18058
rect 17726 17305 17740 18055
rect 17720 17302 17746 17305
rect 17720 17273 17746 17276
rect 17858 17302 17884 17305
rect 17956 17296 17970 18361
rect 18002 17339 18016 20877
rect 18364 20090 18390 20093
rect 18364 20061 18390 20064
rect 18370 20025 18384 20061
rect 18364 20022 18390 20025
rect 18364 19993 18390 19996
rect 17996 17336 18022 17339
rect 17996 17307 18022 17310
rect 17884 17282 17970 17296
rect 17858 17273 17884 17276
rect 17674 17268 17700 17271
rect 17674 17239 17700 17242
rect 17726 16761 17740 17273
rect 17720 16758 17746 16761
rect 17720 16729 17746 16732
rect 17904 16758 17930 16761
rect 17956 16752 17970 17282
rect 17930 16738 17970 16752
rect 17904 16729 17930 16732
rect 18318 15636 18344 15639
rect 18318 15607 18344 15610
rect 18324 15571 18338 15607
rect 18318 15568 18344 15571
rect 18318 15539 18344 15542
rect 18324 15401 18338 15539
rect 18318 15398 18344 15401
rect 18318 15369 18344 15372
rect 17904 14310 17930 14313
rect 17904 14281 17930 14284
rect 17674 14276 17700 14279
rect 17674 14247 17700 14250
rect 17680 14041 17694 14247
rect 17766 14242 17792 14245
rect 17766 14213 17792 14216
rect 17720 14208 17746 14211
rect 17720 14179 17746 14182
rect 17674 14038 17700 14041
rect 17674 14009 17700 14012
rect 17444 12984 17470 12987
rect 17444 12955 17470 12958
rect 17220 12409 17280 12417
rect 17680 12409 17694 14009
rect 17726 13531 17740 14179
rect 17772 14109 17786 14213
rect 17812 14208 17838 14211
rect 17812 14179 17838 14182
rect 17766 14106 17792 14109
rect 17766 14077 17792 14080
rect 17818 13735 17832 14179
rect 17812 13732 17838 13735
rect 17812 13703 17838 13706
rect 17720 13528 17746 13531
rect 17720 13499 17746 13502
rect 17858 13528 17884 13531
rect 17858 13499 17884 13502
rect 17864 12409 17878 13499
rect 17910 12409 17924 14281
rect 18317 13512 18345 13516
rect 18317 13479 18318 13484
rect 18344 13479 18345 13484
rect 18318 13465 18344 13468
rect 18324 12579 18338 13465
rect 18318 12576 18344 12579
rect 18318 12547 18344 12550
rect 18324 12443 18338 12547
rect 18318 12440 18344 12443
rect 18318 12411 18344 12414
rect 17030 12406 17056 12409
rect 17030 12377 17056 12380
rect 17168 12406 17194 12409
rect 17168 12377 17194 12380
rect 17214 12406 17280 12409
rect 17240 12403 17280 12406
rect 17214 12377 17240 12380
rect 16984 12304 17010 12307
rect 16984 12275 17010 12278
rect 16990 12103 17004 12275
rect 16984 12100 17010 12103
rect 16984 12071 17010 12074
rect 17036 11083 17050 12377
rect 17214 12338 17240 12341
rect 17214 12309 17240 12312
rect 17168 12032 17194 12035
rect 17168 12003 17194 12006
rect 17122 11318 17148 11321
rect 17122 11289 17148 11292
rect 17076 11284 17102 11287
rect 17076 11255 17102 11258
rect 17030 11080 17056 11083
rect 17030 11051 17056 11054
rect 17082 10388 17096 11255
rect 17128 11083 17142 11289
rect 17122 11080 17148 11083
rect 17122 11051 17148 11054
rect 17174 11047 17188 12003
rect 17220 11287 17234 12309
rect 17266 12103 17280 12403
rect 17674 12406 17700 12409
rect 17674 12377 17700 12380
rect 17858 12406 17884 12409
rect 17858 12377 17884 12380
rect 17904 12406 17930 12409
rect 17904 12377 17930 12380
rect 17536 12304 17562 12307
rect 17536 12275 17562 12278
rect 17542 12103 17556 12275
rect 17910 12103 17924 12377
rect 18324 12341 18338 12411
rect 18318 12338 18344 12341
rect 18318 12309 18344 12312
rect 17260 12100 17286 12103
rect 17260 12071 17286 12074
rect 17536 12100 17562 12103
rect 17536 12071 17562 12074
rect 17904 12100 17930 12103
rect 17904 12071 17930 12074
rect 17444 11590 17470 11593
rect 17444 11561 17470 11564
rect 17450 11321 17464 11561
rect 17444 11318 17470 11321
rect 17444 11289 17470 11292
rect 17536 11318 17562 11321
rect 17536 11289 17562 11292
rect 17214 11284 17240 11287
rect 17214 11255 17240 11258
rect 17220 11125 17234 11255
rect 17220 11111 17280 11125
rect 17214 11047 17240 11049
rect 17174 11046 17240 11047
rect 17174 11033 17214 11046
rect 17214 11017 17240 11020
rect 17168 11012 17194 11015
rect 17168 10983 17194 10986
rect 17122 10400 17148 10403
rect 17075 10384 17103 10388
rect 17122 10371 17148 10374
rect 17075 10351 17103 10356
rect 17128 9927 17142 10371
rect 17122 9924 17148 9927
rect 17122 9895 17148 9898
rect 17030 9720 17056 9723
rect 17030 9691 17056 9694
rect 16570 9652 16596 9655
rect 16938 9652 16964 9655
rect 16570 9623 16596 9626
rect 16707 9636 16735 9640
rect 16110 9380 16136 9383
rect 16110 9351 16136 9354
rect 15978 9207 16038 9221
rect 15926 9176 15952 9179
rect 15926 9147 15952 9150
rect 15880 8020 15906 8023
rect 15880 7991 15906 7994
rect 15788 7578 15814 7581
rect 15788 7549 15814 7552
rect 15742 7510 15768 7513
rect 15742 7481 15768 7484
rect 15748 7003 15762 7481
rect 15788 7204 15814 7207
rect 15788 7175 15814 7178
rect 15742 7000 15768 7003
rect 15742 6971 15768 6974
rect 15748 6935 15762 6971
rect 15794 6969 15808 7175
rect 15788 6966 15814 6969
rect 15788 6937 15814 6940
rect 15742 6932 15768 6935
rect 15742 6903 15768 6906
rect 15932 6459 15946 9147
rect 15972 9142 15998 9145
rect 15972 9113 15998 9116
rect 15978 8941 15992 9113
rect 16024 9043 16038 9207
rect 16018 9040 16044 9043
rect 16018 9011 16044 9014
rect 15972 8938 15998 8941
rect 15972 8909 15998 8912
rect 16576 8805 16590 9623
rect 16938 9623 16964 9626
rect 16707 9603 16735 9608
rect 16570 8802 16596 8805
rect 16570 8773 16596 8776
rect 16110 8054 16136 8057
rect 16110 8025 16136 8028
rect 15972 8020 15998 8023
rect 15972 7991 15998 7994
rect 15978 7853 15992 7991
rect 15972 7850 15998 7853
rect 15972 7821 15998 7824
rect 15972 7748 15998 7751
rect 15972 7719 15998 7722
rect 15926 6456 15952 6459
rect 15926 6427 15952 6430
rect 15978 6425 15992 7719
rect 16116 6629 16130 8025
rect 16294 6966 16320 6969
rect 16294 6937 16320 6940
rect 16110 6626 16136 6629
rect 16110 6597 16136 6600
rect 16018 6456 16044 6459
rect 16018 6427 16044 6430
rect 15972 6422 15998 6425
rect 15972 6393 15998 6396
rect 15702 6203 15762 6217
rect 15236 5538 15262 5541
rect 15236 5509 15262 5512
rect 15696 5504 15722 5507
rect 15696 5475 15722 5478
rect 15702 5371 15716 5475
rect 15696 5368 15722 5371
rect 15696 5339 15722 5342
rect 13908 3443 13968 3457
rect 13908 0 13922 3443
rect 15748 0 15762 6203
rect 15926 5776 15952 5779
rect 15926 5747 15952 5750
rect 15932 5337 15946 5747
rect 15978 5405 15992 6393
rect 15972 5402 15998 5405
rect 15972 5373 15998 5376
rect 15926 5334 15952 5337
rect 15926 5305 15952 5308
rect 15932 4827 15946 5305
rect 15978 4861 15992 5373
rect 16024 5303 16038 6427
rect 16116 6425 16130 6597
rect 16110 6422 16136 6425
rect 16110 6393 16136 6396
rect 16064 5606 16090 5609
rect 16064 5577 16090 5580
rect 16070 5405 16084 5577
rect 16064 5402 16090 5405
rect 16064 5373 16090 5376
rect 16116 5337 16130 6393
rect 16300 6391 16314 6937
rect 16576 6935 16590 8773
rect 16570 6932 16596 6935
rect 16570 6903 16596 6906
rect 16294 6388 16320 6391
rect 16294 6359 16320 6362
rect 16524 6320 16550 6323
rect 16524 6291 16550 6294
rect 16530 5609 16544 6291
rect 16576 5643 16590 6903
rect 16570 5640 16596 5643
rect 16570 5611 16596 5614
rect 16524 5606 16550 5609
rect 16524 5577 16550 5580
rect 16110 5334 16136 5337
rect 16110 5305 16136 5308
rect 16018 5300 16044 5303
rect 16018 5271 16044 5274
rect 16024 5235 16038 5271
rect 16018 5232 16044 5235
rect 16018 5203 16044 5206
rect 15972 4858 15998 4861
rect 15972 4829 15998 4832
rect 15926 4824 15952 4827
rect 15926 4795 15952 4798
rect 16714 679 16728 9603
rect 17036 6391 17050 9691
rect 17128 9689 17142 9895
rect 17122 9686 17148 9689
rect 17122 9657 17148 9660
rect 17128 9111 17142 9657
rect 17174 9111 17188 10983
rect 17266 10981 17280 11111
rect 17260 10978 17286 10981
rect 17260 10949 17286 10952
rect 17266 10573 17280 10949
rect 17542 10743 17556 11289
rect 17904 11012 17930 11015
rect 17904 10983 17930 10986
rect 17536 10740 17562 10743
rect 17536 10711 17562 10714
rect 17260 10570 17286 10573
rect 17260 10541 17286 10544
rect 17214 10468 17240 10471
rect 17214 10439 17240 10442
rect 17220 10199 17234 10439
rect 17214 10196 17240 10199
rect 17214 10167 17240 10170
rect 17220 9927 17234 10167
rect 17910 9961 17924 10983
rect 18324 10981 18338 12309
rect 18318 10978 18344 10981
rect 18318 10949 18344 10952
rect 18324 10743 18338 10949
rect 18318 10740 18344 10743
rect 18318 10711 18344 10714
rect 18324 9961 18338 10711
rect 17904 9958 17930 9961
rect 17904 9929 17930 9932
rect 18318 9958 18344 9961
rect 18318 9929 18344 9932
rect 17214 9924 17240 9927
rect 17214 9895 17240 9898
rect 17858 9924 17884 9927
rect 17858 9895 17884 9898
rect 17220 9723 17234 9895
rect 17214 9720 17240 9723
rect 17214 9691 17240 9694
rect 17076 9108 17102 9111
rect 17076 9079 17102 9082
rect 17122 9108 17148 9111
rect 17122 9079 17148 9082
rect 17168 9108 17194 9111
rect 17168 9079 17194 9082
rect 17082 8805 17096 9079
rect 17076 8802 17102 8805
rect 17076 8773 17102 8776
rect 17082 8601 17096 8773
rect 17128 8745 17142 9079
rect 17168 9040 17194 9043
rect 17168 9011 17194 9014
rect 17174 8839 17188 9011
rect 17864 8941 17878 9895
rect 17858 8938 17884 8941
rect 17858 8909 17884 8912
rect 18226 8870 18252 8873
rect 18226 8841 18252 8844
rect 17168 8836 17194 8839
rect 17168 8807 17194 8810
rect 17996 8836 18022 8839
rect 17996 8807 18022 8810
rect 17128 8731 17188 8745
rect 17174 8601 17188 8731
rect 17076 8598 17102 8601
rect 17076 8569 17102 8572
rect 17168 8598 17194 8601
rect 17168 8569 17194 8572
rect 17122 8530 17148 8533
rect 17122 8501 17148 8504
rect 17128 6425 17142 8501
rect 17174 7989 17188 8569
rect 18002 8125 18016 8807
rect 18232 8601 18246 8841
rect 18226 8598 18252 8601
rect 18226 8569 18252 8572
rect 18272 8564 18298 8567
rect 18272 8535 18298 8538
rect 18278 8125 18292 8535
rect 18370 8287 18384 19993
rect 18416 15129 18430 23019
rect 18554 23017 18568 23529
rect 18600 23493 18614 23971
rect 19376 23830 19402 23833
rect 19376 23801 19402 23804
rect 19382 23561 19396 23801
rect 19376 23558 19402 23561
rect 19376 23529 19402 23532
rect 18594 23490 18620 23493
rect 18594 23461 18620 23464
rect 18548 23014 18574 23017
rect 18548 22985 18574 22988
rect 18554 22779 18568 22985
rect 18548 22776 18574 22779
rect 18548 22747 18574 22750
rect 18600 22702 18614 23461
rect 19382 23221 19396 23529
rect 19428 23493 19442 24617
rect 19422 23490 19448 23493
rect 19422 23461 19448 23464
rect 19428 23289 19442 23461
rect 19422 23286 19448 23289
rect 19422 23257 19448 23260
rect 19376 23218 19402 23221
rect 19376 23189 19402 23192
rect 18640 22708 18666 22711
rect 18584 22688 18640 22702
rect 18584 22685 18598 22688
rect 18508 22671 18598 22685
rect 18640 22679 18666 22682
rect 18508 22643 18522 22671
rect 18584 22668 18598 22671
rect 19192 22674 19218 22677
rect 18584 22654 18614 22668
rect 18502 22640 18528 22643
rect 18502 22611 18528 22614
rect 18548 22640 18574 22643
rect 18548 22611 18574 22614
rect 18502 22402 18528 22405
rect 18502 22373 18528 22376
rect 18508 22133 18522 22373
rect 18554 22235 18568 22611
rect 18600 22269 18614 22654
rect 19192 22645 19218 22648
rect 18594 22266 18620 22269
rect 18594 22237 18620 22240
rect 18548 22232 18574 22235
rect 18548 22203 18574 22206
rect 18502 22130 18528 22133
rect 18502 22101 18528 22104
rect 18548 21144 18574 21147
rect 18548 21115 18574 21118
rect 18554 20909 18568 21115
rect 19008 21008 19034 21011
rect 19008 20979 19034 20982
rect 18548 20906 18574 20909
rect 18548 20877 18574 20880
rect 19014 20841 19028 20979
rect 19008 20838 19034 20841
rect 19008 20809 19034 20812
rect 18870 19920 18896 19923
rect 18870 19891 18896 19894
rect 18640 19172 18666 19175
rect 18640 19143 18666 19146
rect 18456 18662 18482 18665
rect 18456 18633 18482 18636
rect 18462 18393 18476 18633
rect 18456 18390 18482 18393
rect 18456 18361 18482 18364
rect 18646 15760 18660 19143
rect 18685 18476 18713 18480
rect 18685 18443 18713 18448
rect 18639 15756 18667 15760
rect 18600 15735 18639 15749
rect 18600 15707 18614 15735
rect 18639 15723 18667 15728
rect 18594 15704 18620 15707
rect 18594 15675 18620 15678
rect 18692 15333 18706 18443
rect 18876 17849 18890 19891
rect 19146 18832 19172 18835
rect 19146 18803 19172 18806
rect 18915 18476 18943 18480
rect 18915 18443 18943 18448
rect 18922 18393 18936 18443
rect 18916 18390 18942 18393
rect 18916 18361 18942 18364
rect 18778 17846 18804 17849
rect 18778 17817 18804 17820
rect 18870 17846 18896 17849
rect 18870 17817 18896 17820
rect 18784 17645 18798 17817
rect 18778 17642 18804 17645
rect 18778 17613 18804 17616
rect 19008 17608 19034 17611
rect 19008 17579 19034 17582
rect 18824 17540 18850 17543
rect 18824 17511 18850 17514
rect 18916 17540 18942 17543
rect 19014 17532 19028 17579
rect 19152 17577 19166 18803
rect 19146 17574 19172 17577
rect 19146 17545 19172 17548
rect 18916 17511 18942 17514
rect 18991 17529 19028 17532
rect 18830 16829 18844 17511
rect 18922 17373 18936 17511
rect 19017 17503 19028 17529
rect 18991 17500 19017 17503
rect 18997 17466 19011 17500
rect 18968 17452 19011 17466
rect 19100 17472 19126 17475
rect 18916 17370 18942 17373
rect 18916 17341 18942 17344
rect 18824 16826 18850 16829
rect 18824 16797 18850 16800
rect 18732 15670 18758 15673
rect 18732 15641 18758 15644
rect 18738 15367 18752 15641
rect 18916 15466 18942 15469
rect 18916 15437 18942 15440
rect 18732 15364 18758 15367
rect 18732 15335 18758 15338
rect 18870 15364 18896 15367
rect 18870 15335 18896 15338
rect 18686 15330 18712 15333
rect 18686 15301 18712 15304
rect 18410 15126 18436 15129
rect 18410 15097 18436 15100
rect 18416 11321 18430 15097
rect 18824 13698 18850 13701
rect 18824 13669 18850 13672
rect 18732 13426 18758 13429
rect 18732 13397 18758 13400
rect 18778 13426 18804 13429
rect 18778 13397 18804 13400
rect 18738 13191 18752 13397
rect 18686 13188 18712 13191
rect 18686 13159 18712 13162
rect 18732 13188 18758 13191
rect 18732 13159 18758 13162
rect 18692 13114 18706 13159
rect 18784 13114 18798 13397
rect 18830 13293 18844 13669
rect 18824 13290 18850 13293
rect 18824 13261 18850 13264
rect 18692 13100 18798 13114
rect 18594 12372 18620 12375
rect 18594 12343 18620 12346
rect 18502 12304 18528 12307
rect 18502 12275 18528 12278
rect 18508 12137 18522 12275
rect 18502 12134 18528 12137
rect 18502 12105 18528 12108
rect 18548 11522 18574 11525
rect 18548 11493 18574 11496
rect 18554 11321 18568 11493
rect 18600 11355 18614 12343
rect 18640 12134 18666 12137
rect 18640 12105 18666 12108
rect 18646 11559 18660 12105
rect 18732 11862 18758 11865
rect 18732 11833 18758 11836
rect 18738 11661 18752 11833
rect 18732 11658 18758 11661
rect 18732 11629 18758 11632
rect 18640 11556 18666 11559
rect 18640 11527 18666 11530
rect 18732 11556 18758 11559
rect 18732 11527 18758 11530
rect 18594 11352 18620 11355
rect 18594 11323 18620 11326
rect 18410 11318 18436 11321
rect 18410 11289 18436 11292
rect 18548 11318 18574 11321
rect 18548 11289 18574 11292
rect 18594 11216 18620 11219
rect 18594 11187 18620 11190
rect 18600 11015 18614 11187
rect 18738 11117 18752 11527
rect 18732 11114 18758 11117
rect 18732 11085 18758 11088
rect 18738 11047 18752 11085
rect 18692 11033 18752 11047
rect 18594 11012 18620 11015
rect 18594 10983 18620 10986
rect 18640 10672 18666 10675
rect 18640 10643 18666 10646
rect 18646 10471 18660 10643
rect 18692 10471 18706 11033
rect 18732 10774 18758 10777
rect 18732 10745 18758 10748
rect 18738 10573 18752 10745
rect 18732 10570 18758 10573
rect 18732 10541 18758 10544
rect 18640 10468 18666 10471
rect 18640 10439 18666 10442
rect 18686 10468 18712 10471
rect 18686 10439 18712 10442
rect 18640 9380 18666 9383
rect 18640 9351 18666 9354
rect 18646 9179 18660 9351
rect 18640 9176 18666 9179
rect 18640 9147 18666 9150
rect 18410 8768 18436 8771
rect 18410 8739 18436 8742
rect 18416 8669 18430 8739
rect 18410 8666 18436 8669
rect 18410 8637 18436 8640
rect 18370 8273 18430 8287
rect 17996 8122 18022 8125
rect 17996 8093 18022 8096
rect 18272 8122 18298 8125
rect 18272 8093 18298 8096
rect 17490 8054 17516 8057
rect 17490 8025 17516 8028
rect 18088 8054 18114 8057
rect 18088 8025 18114 8028
rect 17398 8020 17424 8023
rect 17398 7991 17424 7994
rect 17168 7986 17194 7989
rect 17168 7957 17194 7960
rect 17404 6901 17418 7991
rect 17496 7853 17510 8025
rect 17490 7850 17516 7853
rect 17490 7821 17516 7824
rect 18094 6969 18108 8025
rect 18272 7782 18298 7785
rect 18272 7753 18298 7756
rect 18278 7581 18292 7753
rect 18318 7748 18344 7751
rect 18318 7719 18344 7722
rect 18272 7578 18298 7581
rect 18272 7549 18298 7552
rect 18324 7513 18338 7719
rect 18318 7510 18344 7513
rect 18318 7481 18344 7484
rect 18324 7249 18338 7481
rect 18324 7235 18384 7249
rect 18318 7170 18344 7173
rect 18318 7141 18344 7144
rect 18324 6969 18338 7141
rect 17858 6966 17884 6969
rect 17858 6937 17884 6940
rect 18088 6966 18114 6969
rect 18088 6937 18114 6940
rect 18318 6966 18344 6969
rect 18318 6937 18344 6940
rect 17398 6898 17424 6901
rect 17398 6869 17424 6872
rect 17864 6663 17878 6937
rect 18094 6663 18108 6937
rect 17858 6660 17884 6663
rect 17858 6631 17884 6634
rect 18088 6660 18114 6663
rect 18088 6631 18114 6634
rect 17864 6459 17878 6631
rect 17858 6456 17884 6459
rect 17858 6427 17884 6430
rect 17122 6422 17148 6425
rect 17122 6393 17148 6396
rect 17030 6388 17056 6391
rect 17030 6359 17056 6362
rect 17036 5881 17050 6359
rect 17128 5881 17142 6393
rect 18094 5915 18108 6631
rect 18134 6592 18160 6595
rect 18134 6563 18160 6566
rect 18140 6425 18154 6563
rect 18134 6422 18160 6425
rect 18134 6393 18160 6396
rect 18088 5912 18114 5915
rect 18088 5883 18114 5886
rect 17030 5878 17056 5881
rect 17030 5849 17056 5852
rect 17122 5878 17148 5881
rect 17122 5849 17148 5852
rect 17214 5878 17240 5881
rect 17214 5849 17240 5852
rect 18272 5878 18298 5881
rect 18272 5849 18298 5852
rect 17030 5606 17056 5609
rect 17030 5577 17056 5580
rect 16984 5504 17010 5507
rect 16984 5475 17010 5478
rect 16990 5337 17004 5475
rect 16984 5334 17010 5337
rect 16984 5305 17010 5308
rect 17036 5269 17050 5577
rect 17122 5538 17148 5541
rect 17122 5509 17148 5512
rect 17128 5371 17142 5509
rect 17122 5368 17148 5371
rect 17122 5339 17148 5342
rect 17030 5266 17056 5269
rect 17030 5237 17056 5240
rect 17036 4793 17050 5237
rect 17030 4790 17056 4793
rect 17030 4761 17056 4764
rect 17128 4759 17142 5339
rect 17220 4793 17234 5849
rect 18278 5541 18292 5849
rect 17398 5538 17424 5541
rect 17398 5509 17424 5512
rect 18272 5538 18298 5541
rect 18272 5509 18298 5512
rect 17404 5405 17418 5509
rect 17398 5402 17424 5405
rect 17398 5373 17424 5376
rect 18278 5337 18292 5509
rect 18272 5334 18298 5337
rect 18272 5305 18298 5308
rect 18278 5065 18292 5305
rect 18318 5300 18344 5303
rect 18318 5271 18344 5274
rect 18370 5277 18384 7235
rect 18416 7139 18430 8273
rect 18646 8057 18660 9147
rect 18640 8054 18666 8057
rect 18640 8025 18666 8028
rect 18646 7207 18660 8025
rect 18640 7204 18666 7207
rect 18640 7175 18666 7178
rect 18410 7136 18436 7139
rect 18410 7107 18436 7110
rect 18410 7000 18436 7003
rect 18410 6971 18436 6974
rect 18416 6425 18430 6971
rect 18876 6935 18890 15335
rect 18922 15129 18936 15437
rect 18916 15126 18942 15129
rect 18916 15097 18942 15100
rect 18968 11047 18982 17452
rect 19100 17443 19126 17446
rect 19053 13512 19081 13516
rect 19053 13479 19054 13484
rect 19080 13479 19081 13484
rect 19054 13465 19080 13468
rect 18922 11033 18982 11047
rect 18922 9111 18936 11033
rect 19106 10241 19120 17443
rect 19146 12406 19172 12409
rect 19146 12377 19172 12380
rect 19152 12205 19166 12377
rect 19146 12202 19172 12205
rect 19146 12173 19172 12176
rect 18968 10227 19120 10241
rect 18968 9315 18982 10227
rect 19054 9992 19080 9995
rect 19054 9963 19080 9966
rect 19008 9652 19034 9655
rect 19008 9623 19034 9626
rect 19014 9417 19028 9623
rect 19008 9414 19034 9417
rect 19008 9385 19034 9388
rect 18962 9312 18988 9315
rect 18962 9283 18988 9286
rect 18916 9108 18942 9111
rect 18916 9079 18942 9082
rect 19060 8805 19074 9963
rect 19100 9686 19126 9689
rect 19100 9657 19126 9660
rect 19146 9686 19172 9689
rect 19146 9657 19172 9660
rect 19106 9383 19120 9657
rect 19100 9380 19126 9383
rect 19100 9351 19126 9354
rect 19152 9349 19166 9657
rect 19146 9346 19172 9349
rect 19146 9317 19172 9320
rect 19152 9145 19166 9317
rect 19146 9142 19172 9145
rect 19146 9113 19172 9116
rect 19054 8802 19080 8805
rect 19054 8773 19080 8776
rect 19100 8258 19126 8261
rect 19100 8229 19126 8232
rect 19106 7717 19120 8229
rect 19146 7748 19172 7751
rect 19146 7719 19172 7722
rect 19100 7714 19126 7717
rect 19100 7685 19126 7688
rect 19106 7513 19120 7685
rect 18962 7510 18988 7513
rect 18962 7481 18988 7484
rect 19100 7510 19126 7513
rect 19100 7481 19126 7484
rect 18968 7241 18982 7481
rect 18962 7238 18988 7241
rect 18962 7209 18988 7212
rect 18870 6932 18896 6935
rect 18870 6903 18896 6906
rect 18968 6663 18982 7209
rect 18962 6660 18988 6663
rect 18962 6631 18988 6634
rect 18410 6422 18436 6425
rect 18410 6393 18436 6396
rect 18416 6217 18430 6393
rect 18686 6388 18712 6391
rect 18686 6359 18712 6362
rect 18416 6203 18522 6217
rect 18508 5881 18522 6203
rect 18548 5946 18574 5949
rect 18548 5917 18574 5920
rect 18502 5878 18528 5881
rect 18502 5849 18528 5852
rect 18508 5575 18522 5849
rect 18554 5575 18568 5917
rect 18692 5677 18706 6359
rect 18686 5674 18712 5677
rect 18686 5645 18712 5648
rect 18502 5572 18528 5575
rect 18502 5543 18528 5546
rect 18548 5572 18574 5575
rect 18548 5543 18574 5546
rect 18968 5337 18982 6631
rect 19106 5915 19120 7481
rect 19152 7241 19166 7719
rect 19146 7238 19172 7241
rect 19146 7209 19172 7212
rect 19152 6663 19166 7209
rect 19146 6660 19172 6663
rect 19146 6631 19172 6634
rect 19152 6459 19166 6631
rect 19146 6456 19172 6459
rect 19146 6427 19172 6430
rect 19100 5912 19126 5915
rect 19100 5883 19126 5886
rect 18962 5334 18988 5337
rect 18962 5305 18988 5308
rect 18272 5062 18298 5065
rect 18272 5033 18298 5036
rect 18324 4861 18338 5271
rect 18370 5263 18476 5277
rect 18462 4963 18476 5263
rect 18640 5232 18666 5235
rect 18640 5203 18666 5206
rect 18646 5031 18660 5203
rect 18968 5065 18982 5305
rect 18962 5062 18988 5065
rect 18962 5033 18988 5036
rect 18640 5028 18666 5031
rect 18640 4999 18666 5002
rect 18456 4960 18482 4963
rect 18456 4931 18482 4934
rect 18594 4960 18620 4963
rect 18594 4931 18620 4934
rect 18318 4858 18344 4861
rect 18318 4829 18344 4832
rect 17260 4824 17286 4827
rect 17260 4795 17286 4798
rect 17214 4790 17240 4793
rect 17214 4761 17240 4764
rect 17122 4756 17148 4759
rect 17122 4727 17148 4730
rect 17076 4688 17102 4691
rect 17076 4659 17102 4662
rect 17082 4487 17096 4659
rect 17128 4589 17142 4727
rect 17266 4589 17280 4795
rect 18462 4793 18476 4931
rect 18600 4827 18614 4931
rect 18594 4824 18620 4827
rect 18594 4795 18620 4798
rect 18456 4790 18482 4793
rect 18456 4761 18482 4764
rect 17122 4586 17148 4589
rect 17122 4557 17148 4560
rect 17260 4586 17286 4589
rect 17260 4557 17286 4560
rect 17076 4484 17102 4487
rect 17076 4455 17102 4458
rect 19198 3977 19212 22645
rect 19382 21929 19396 23189
rect 19376 21926 19402 21929
rect 19376 21897 19402 21900
rect 19382 21869 19396 21897
rect 19336 21855 19396 21869
rect 19336 21385 19350 21855
rect 19474 21589 19488 25523
rect 20256 24615 20270 26011
rect 20486 26009 20500 29063
rect 20900 28805 20914 33000
rect 20900 28797 20960 28805
rect 20900 28794 20966 28797
rect 20900 28791 20940 28794
rect 20848 28726 20874 28729
rect 20848 28697 20874 28700
rect 20618 28454 20644 28457
rect 20618 28425 20644 28428
rect 20526 28352 20552 28355
rect 20526 28323 20552 28326
rect 20532 26213 20546 28323
rect 20624 27913 20638 28425
rect 20854 28219 20868 28697
rect 20900 28423 20914 28791
rect 20940 28765 20966 28768
rect 20894 28420 20920 28423
rect 20894 28391 20920 28394
rect 20710 28216 20736 28219
rect 20710 28187 20736 28190
rect 20848 28216 20874 28219
rect 20848 28187 20874 28190
rect 20618 27910 20644 27913
rect 20618 27881 20644 27884
rect 20572 27808 20598 27811
rect 20572 27779 20598 27782
rect 20578 27437 20592 27779
rect 20624 27607 20638 27881
rect 20624 27593 20684 27607
rect 20572 27434 20598 27437
rect 20572 27405 20598 27408
rect 20618 26720 20644 26723
rect 20618 26691 20644 26694
rect 20624 26621 20638 26691
rect 20618 26618 20644 26621
rect 20618 26589 20644 26592
rect 20670 26519 20684 27593
rect 20716 27131 20730 28187
rect 20992 27607 21006 33000
rect 21084 28253 21098 33000
rect 21078 28250 21104 28253
rect 21078 28221 21104 28224
rect 21084 27879 21098 28221
rect 21078 27876 21104 27879
rect 21078 27847 21104 27850
rect 20992 27593 21144 27607
rect 20710 27128 20736 27131
rect 20710 27099 20736 27102
rect 21130 27063 21144 27593
rect 21308 27128 21334 27131
rect 21308 27099 21334 27102
rect 21124 27060 21150 27063
rect 21124 27031 21150 27034
rect 21130 26587 21144 27031
rect 21124 26584 21150 26587
rect 21124 26555 21150 26558
rect 20664 26516 20690 26519
rect 20664 26487 20690 26490
rect 20526 26210 20552 26213
rect 20526 26181 20552 26184
rect 20480 26006 20506 26009
rect 20480 25977 20506 25980
rect 20486 25703 20500 25977
rect 21078 25972 21104 25975
rect 21078 25943 21104 25946
rect 20480 25700 20506 25703
rect 20480 25671 20506 25674
rect 20486 25159 20500 25671
rect 20480 25156 20506 25159
rect 20480 25127 20506 25130
rect 20388 25088 20414 25091
rect 20388 25059 20414 25062
rect 20394 24887 20408 25059
rect 20388 24884 20414 24887
rect 20388 24855 20414 24858
rect 20342 24816 20368 24819
rect 20342 24787 20368 24790
rect 19560 24612 19586 24615
rect 19560 24583 19586 24586
rect 20250 24612 20276 24615
rect 20250 24583 20276 24586
rect 19566 23833 19580 24583
rect 19606 24578 19632 24581
rect 19606 24549 19632 24552
rect 19612 24377 19626 24549
rect 19606 24374 19632 24377
rect 19606 24345 19632 24348
rect 19560 23830 19586 23833
rect 19560 23801 19586 23804
rect 19612 22745 19626 24345
rect 20020 24068 20046 24071
rect 20020 24039 20046 24042
rect 20026 23527 20040 24039
rect 20020 23524 20046 23527
rect 20020 23495 20046 23498
rect 19652 23014 19678 23017
rect 19652 22985 19678 22988
rect 19658 22813 19672 22985
rect 19790 22946 19816 22949
rect 19790 22917 19816 22920
rect 19652 22810 19678 22813
rect 19652 22781 19678 22784
rect 19606 22742 19632 22745
rect 19606 22713 19632 22716
rect 19796 21895 19810 22917
rect 19790 21892 19816 21895
rect 19790 21863 19816 21866
rect 19468 21586 19494 21589
rect 19468 21557 19494 21560
rect 19330 21382 19356 21385
rect 19330 21353 19356 21356
rect 19284 21314 19310 21317
rect 19284 21285 19310 21288
rect 19290 21079 19304 21285
rect 19284 21076 19310 21079
rect 19284 21047 19310 21050
rect 19238 21042 19264 21045
rect 19238 21013 19264 21016
rect 19244 20773 19258 21013
rect 19290 20807 19304 21047
rect 19336 21011 19350 21353
rect 19560 21314 19586 21317
rect 19560 21285 19586 21288
rect 19330 21008 19356 21011
rect 19330 20979 19356 20982
rect 19284 20804 19310 20807
rect 19284 20775 19310 20778
rect 19238 20770 19264 20773
rect 19238 20741 19264 20744
rect 19244 20093 19258 20741
rect 19336 20297 19350 20979
rect 19376 20362 19402 20365
rect 19376 20333 19402 20336
rect 19330 20294 19356 20297
rect 19330 20265 19356 20268
rect 19238 20090 19264 20093
rect 19238 20061 19264 20064
rect 19336 19753 19350 20265
rect 19382 20229 19396 20333
rect 19566 20263 19580 21285
rect 19796 20365 19810 21863
rect 19790 20362 19816 20365
rect 19790 20333 19816 20336
rect 19560 20260 19586 20263
rect 19560 20231 19586 20234
rect 19376 20226 19402 20229
rect 19376 20197 19402 20200
rect 19330 19750 19356 19753
rect 19330 19721 19356 19724
rect 19336 19277 19350 19721
rect 19382 19685 19396 20197
rect 19376 19682 19402 19685
rect 19376 19653 19402 19656
rect 19238 19274 19264 19277
rect 19238 19245 19264 19248
rect 19330 19274 19356 19277
rect 19330 19245 19356 19248
rect 19244 18631 19258 19245
rect 19382 18631 19396 19653
rect 19238 18628 19264 18631
rect 19238 18599 19264 18602
rect 19376 18628 19402 18631
rect 19376 18599 19402 18602
rect 19244 18291 19258 18599
rect 19238 18288 19264 18291
rect 19238 18259 19264 18262
rect 19382 18019 19396 18599
rect 19376 18016 19402 18019
rect 19376 17987 19402 17990
rect 19284 17744 19310 17747
rect 19284 17715 19310 17718
rect 19290 14313 19304 17715
rect 19928 17540 19954 17543
rect 19928 17511 19954 17514
rect 19652 17302 19678 17305
rect 19652 17273 19678 17276
rect 19284 14310 19310 14313
rect 19284 14281 19310 14284
rect 19376 14276 19402 14279
rect 19376 14247 19402 14250
rect 19382 14075 19396 14247
rect 19514 14208 19540 14211
rect 19514 14179 19540 14182
rect 19376 14072 19402 14075
rect 19376 14043 19402 14046
rect 19382 13667 19396 14043
rect 19376 13664 19402 13667
rect 19376 13635 19402 13638
rect 19382 13565 19396 13635
rect 19376 13562 19402 13565
rect 19376 13533 19402 13536
rect 19520 13531 19534 14179
rect 19514 13528 19540 13531
rect 19514 13499 19540 13502
rect 19284 13154 19310 13157
rect 19284 13125 19310 13128
rect 19290 13021 19304 13125
rect 19284 13018 19310 13021
rect 19284 12989 19310 12992
rect 19238 12984 19264 12987
rect 19237 12968 19238 12972
rect 19264 12968 19265 12972
rect 19237 12935 19265 12940
rect 19376 12950 19402 12953
rect 19376 12921 19402 12924
rect 19284 12916 19310 12919
rect 19284 12887 19310 12890
rect 19290 12171 19304 12887
rect 19382 12341 19396 12921
rect 19514 12644 19540 12647
rect 19514 12615 19540 12618
rect 19376 12338 19402 12341
rect 19376 12309 19402 12312
rect 19422 12304 19448 12307
rect 19422 12275 19448 12278
rect 19284 12168 19310 12171
rect 19284 12139 19310 12142
rect 19376 12066 19402 12069
rect 19428 12060 19442 12275
rect 19520 12171 19534 12615
rect 19514 12168 19540 12171
rect 19514 12139 19540 12142
rect 19402 12046 19442 12060
rect 19376 12037 19402 12040
rect 19382 11933 19396 12037
rect 19468 12032 19494 12035
rect 19468 12003 19494 12006
rect 19376 11930 19402 11933
rect 19376 11901 19402 11904
rect 19474 11559 19488 12003
rect 19468 11556 19494 11559
rect 19468 11527 19494 11530
rect 19330 10672 19356 10675
rect 19330 10643 19356 10646
rect 19336 10505 19350 10643
rect 19330 10502 19356 10505
rect 19330 10473 19356 10476
rect 19336 9927 19350 10473
rect 19658 10437 19672 17273
rect 19882 14276 19908 14279
rect 19882 14247 19908 14250
rect 19888 14109 19902 14247
rect 19882 14106 19908 14109
rect 19882 14077 19908 14080
rect 19888 14041 19902 14077
rect 19882 14038 19908 14041
rect 19882 14009 19908 14012
rect 19888 12681 19902 14009
rect 19882 12678 19908 12681
rect 19882 12649 19908 12652
rect 19888 12145 19902 12649
rect 19842 12131 19902 12145
rect 19842 11559 19856 12131
rect 19882 12100 19908 12103
rect 19882 12071 19908 12074
rect 19836 11556 19862 11559
rect 19836 11527 19862 11530
rect 19652 10434 19678 10437
rect 19652 10405 19678 10408
rect 19330 9924 19356 9927
rect 19330 9895 19356 9898
rect 19238 9720 19264 9723
rect 19238 9691 19264 9694
rect 19244 9213 19258 9691
rect 19336 9667 19350 9895
rect 19336 9653 19396 9667
rect 19284 9380 19310 9383
rect 19284 9351 19310 9354
rect 19238 9210 19264 9213
rect 19238 9181 19264 9184
rect 19238 9142 19264 9145
rect 19238 9113 19264 9116
rect 19244 8601 19258 9113
rect 19290 9077 19304 9351
rect 19382 9111 19396 9653
rect 19606 9380 19632 9383
rect 19606 9351 19632 9354
rect 19612 9145 19626 9351
rect 19606 9142 19632 9145
rect 19606 9113 19632 9116
rect 19376 9108 19402 9111
rect 19376 9079 19402 9082
rect 19284 9074 19310 9077
rect 19284 9045 19310 9048
rect 19238 8598 19264 8601
rect 19238 8569 19264 8572
rect 19244 8363 19258 8569
rect 19238 8360 19264 8363
rect 19238 8331 19264 8334
rect 19290 8125 19304 9045
rect 19606 8292 19632 8295
rect 19606 8263 19632 8266
rect 19284 8122 19310 8125
rect 19284 8093 19310 8096
rect 19290 7819 19304 8093
rect 19330 8020 19356 8023
rect 19330 7991 19356 7994
rect 19284 7816 19310 7819
rect 19284 7787 19310 7790
rect 19336 7513 19350 7991
rect 19330 7510 19356 7513
rect 19330 7481 19356 7484
rect 19336 6663 19350 7481
rect 19612 7207 19626 8263
rect 19658 7853 19672 10405
rect 19888 9621 19902 12071
rect 19934 11763 19948 17511
rect 19974 15568 20000 15571
rect 19974 15539 20000 15542
rect 19980 15333 19994 15539
rect 19974 15330 20000 15333
rect 19974 15301 20000 15304
rect 19974 14038 20000 14041
rect 19974 14009 20000 14012
rect 19980 12647 19994 14009
rect 19974 12644 20000 12647
rect 19974 12615 20000 12618
rect 19928 11760 19954 11763
rect 19928 11731 19954 11734
rect 19928 11556 19954 11559
rect 19928 11527 19954 11530
rect 19934 10811 19948 11527
rect 19928 10808 19954 10811
rect 19928 10779 19954 10782
rect 19934 10709 19948 10779
rect 19928 10706 19954 10709
rect 19928 10677 19954 10680
rect 20026 10403 20040 23495
rect 20348 22983 20362 24787
rect 20388 24544 20414 24547
rect 20388 24515 20414 24518
rect 20394 24343 20408 24515
rect 21084 24445 21098 25943
rect 21078 24442 21104 24445
rect 21078 24413 21104 24416
rect 20986 24374 21012 24377
rect 20986 24345 21012 24348
rect 20388 24340 20414 24343
rect 20388 24311 20414 24314
rect 20992 24139 21006 24345
rect 21170 24340 21196 24343
rect 21170 24311 21196 24314
rect 20986 24136 21012 24139
rect 20986 24107 21012 24110
rect 20434 24102 20460 24105
rect 20434 24073 20460 24076
rect 20440 23629 20454 24073
rect 20434 23626 20460 23629
rect 20434 23597 20460 23600
rect 21078 23286 21104 23289
rect 21078 23257 21104 23260
rect 21084 23051 21098 23257
rect 21124 23184 21150 23187
rect 21124 23155 21150 23158
rect 21078 23048 21104 23051
rect 21078 23019 21104 23022
rect 21130 22983 21144 23155
rect 20158 22980 20184 22983
rect 20158 22951 20184 22954
rect 20342 22980 20368 22983
rect 20342 22951 20368 22954
rect 21124 22980 21150 22983
rect 21124 22951 21150 22954
rect 20164 22677 20178 22951
rect 20848 22912 20874 22915
rect 20848 22883 20874 22886
rect 20158 22674 20184 22677
rect 20158 22645 20184 22648
rect 20664 21824 20690 21827
rect 20664 21795 20690 21798
rect 20388 21416 20414 21419
rect 20388 21387 20414 21390
rect 20342 21348 20368 21351
rect 20342 21319 20368 21322
rect 20112 21280 20138 21283
rect 20112 21251 20138 21254
rect 20118 21113 20132 21251
rect 20348 21147 20362 21319
rect 20394 21181 20408 21387
rect 20388 21178 20414 21181
rect 20388 21149 20414 21152
rect 20342 21144 20368 21147
rect 20480 21144 20506 21147
rect 20342 21115 20368 21118
rect 20394 21118 20480 21121
rect 20394 21115 20506 21118
rect 20112 21110 20138 21113
rect 20112 21081 20138 21084
rect 20250 21110 20276 21113
rect 20250 21081 20276 21084
rect 20066 19512 20092 19515
rect 20066 19483 20092 19486
rect 20072 15469 20086 19483
rect 20118 17611 20132 21081
rect 20256 20909 20270 21081
rect 20250 20906 20276 20909
rect 20250 20877 20276 20880
rect 20348 20025 20362 21115
rect 20394 21107 20500 21115
rect 20394 21045 20408 21107
rect 20388 21042 20414 21045
rect 20388 21013 20414 21016
rect 20434 21042 20460 21045
rect 20434 21013 20460 21016
rect 20440 20875 20454 21013
rect 20434 20872 20460 20875
rect 20434 20843 20460 20846
rect 20670 20025 20684 21795
rect 20802 20192 20828 20195
rect 20802 20163 20828 20166
rect 20808 20059 20822 20163
rect 20802 20056 20828 20059
rect 20802 20027 20828 20030
rect 20342 20022 20368 20025
rect 20342 19993 20368 19996
rect 20572 20022 20598 20025
rect 20572 19993 20598 19996
rect 20664 20022 20690 20025
rect 20664 19993 20690 19996
rect 20756 20022 20782 20025
rect 20756 19993 20782 19996
rect 20434 19648 20460 19651
rect 20434 19619 20460 19622
rect 20440 19515 20454 19619
rect 20578 19549 20592 19993
rect 20762 19976 20776 19993
rect 20755 19972 20783 19976
rect 20755 19939 20783 19944
rect 20664 19920 20690 19923
rect 20664 19891 20690 19894
rect 20572 19546 20598 19549
rect 20572 19517 20598 19520
rect 20434 19512 20460 19515
rect 20434 19483 20460 19486
rect 20296 19478 20322 19481
rect 20296 19449 20322 19452
rect 20302 19277 20316 19449
rect 20296 19274 20322 19277
rect 20296 19245 20322 19248
rect 20670 18665 20684 19891
rect 20710 19206 20736 19209
rect 20710 19177 20736 19180
rect 20716 18937 20730 19177
rect 20710 18934 20736 18937
rect 20710 18905 20736 18908
rect 20664 18662 20690 18665
rect 20664 18633 20690 18636
rect 20480 18628 20506 18631
rect 20506 18608 20546 18622
rect 20480 18599 20506 18602
rect 20341 18544 20369 18548
rect 20341 18511 20369 18516
rect 20158 18016 20184 18019
rect 20158 17987 20184 17990
rect 20164 17849 20178 17987
rect 20158 17846 20184 17849
rect 20158 17817 20184 17820
rect 20112 17608 20138 17611
rect 20112 17579 20138 17582
rect 20164 17305 20178 17817
rect 20158 17302 20184 17305
rect 20158 17273 20184 17276
rect 20111 16912 20139 16916
rect 20111 16879 20139 16884
rect 20118 16772 20132 16879
rect 20112 16769 20138 16772
rect 20164 16761 20178 17273
rect 20112 16740 20138 16743
rect 20158 16758 20184 16761
rect 20118 15707 20132 16740
rect 20158 16729 20184 16732
rect 20112 15704 20138 15707
rect 20112 15675 20138 15678
rect 20296 15704 20322 15707
rect 20296 15675 20322 15678
rect 20302 15571 20316 15675
rect 20250 15568 20276 15571
rect 20250 15539 20276 15542
rect 20296 15568 20322 15571
rect 20296 15539 20322 15542
rect 20066 15466 20092 15469
rect 20066 15437 20092 15440
rect 20072 15333 20086 15437
rect 20204 15432 20230 15435
rect 20204 15403 20230 15406
rect 20210 15333 20224 15403
rect 20066 15330 20092 15333
rect 20066 15301 20092 15304
rect 20204 15330 20230 15333
rect 20204 15301 20230 15304
rect 20066 14004 20092 14007
rect 20066 13975 20092 13978
rect 20072 13939 20086 13975
rect 20066 13936 20092 13939
rect 20066 13907 20092 13910
rect 20072 13463 20086 13907
rect 20066 13460 20092 13463
rect 20066 13431 20092 13434
rect 20112 11862 20138 11865
rect 20112 11833 20138 11836
rect 20118 11321 20132 11833
rect 20158 11828 20184 11831
rect 20158 11799 20184 11802
rect 20112 11318 20138 11321
rect 20112 11289 20138 11292
rect 20118 10743 20132 11289
rect 20164 11287 20178 11799
rect 20158 11284 20184 11287
rect 20158 11255 20184 11258
rect 20112 10740 20138 10743
rect 20112 10711 20138 10714
rect 20118 10471 20132 10711
rect 20164 10675 20178 11255
rect 20158 10672 20184 10675
rect 20158 10643 20184 10646
rect 20112 10468 20138 10471
rect 20112 10439 20138 10442
rect 20020 10400 20046 10403
rect 20020 10371 20046 10374
rect 19882 9618 19908 9621
rect 19882 9589 19908 9592
rect 19698 9108 19724 9111
rect 19698 9079 19724 9082
rect 19704 8873 19718 9079
rect 19928 8938 19954 8941
rect 19928 8909 19954 8912
rect 19698 8870 19724 8873
rect 19698 8841 19724 8844
rect 19934 8805 19948 8909
rect 19928 8802 19954 8805
rect 19928 8773 19954 8776
rect 19790 8292 19816 8295
rect 19790 8263 19816 8266
rect 19652 7850 19678 7853
rect 19652 7821 19678 7824
rect 19658 7547 19672 7821
rect 19652 7544 19678 7547
rect 19652 7515 19678 7518
rect 19796 7207 19810 8263
rect 19934 7683 19948 8773
rect 20026 8329 20040 10371
rect 20066 9176 20092 9179
rect 20066 9147 20092 9150
rect 20020 8326 20046 8329
rect 20020 8297 20046 8300
rect 20020 7816 20046 7819
rect 20020 7787 20046 7790
rect 20026 7751 20040 7787
rect 20020 7748 20046 7751
rect 20020 7719 20046 7722
rect 19928 7680 19954 7683
rect 19928 7651 19954 7654
rect 20072 7241 20086 9147
rect 20118 9145 20132 10439
rect 20112 9142 20138 9145
rect 20112 9113 20138 9116
rect 20118 8839 20132 9113
rect 20112 8836 20138 8839
rect 20138 8816 20178 8830
rect 20112 8807 20138 8810
rect 20066 7238 20092 7241
rect 20066 7209 20092 7212
rect 19606 7204 19632 7207
rect 19606 7175 19632 7178
rect 19790 7204 19816 7207
rect 19790 7175 19816 7178
rect 19974 7204 20000 7207
rect 19974 7175 20000 7178
rect 19376 7136 19402 7139
rect 19376 7107 19402 7110
rect 19382 6935 19396 7107
rect 19612 6969 19626 7175
rect 19606 6966 19632 6969
rect 19606 6937 19632 6940
rect 19882 6966 19908 6969
rect 19882 6937 19908 6940
rect 19376 6932 19402 6935
rect 19376 6903 19402 6906
rect 19330 6660 19356 6663
rect 19330 6631 19356 6634
rect 19336 6459 19350 6631
rect 19382 6459 19396 6903
rect 19330 6456 19356 6459
rect 19330 6427 19356 6430
rect 19376 6456 19402 6459
rect 19376 6427 19402 6430
rect 19336 5881 19350 6427
rect 19888 6119 19902 6937
rect 19980 6935 19994 7175
rect 20164 7003 20178 8816
rect 20210 8227 20224 15301
rect 20256 15129 20270 15539
rect 20250 15126 20276 15129
rect 20250 15097 20276 15100
rect 20348 11047 20362 18511
rect 20532 18189 20546 18608
rect 20618 18594 20644 18597
rect 20618 18565 20644 18568
rect 20664 18594 20690 18597
rect 20664 18565 20690 18568
rect 20624 18548 20638 18565
rect 20617 18544 20645 18548
rect 20617 18511 20645 18516
rect 20670 18461 20684 18565
rect 20664 18458 20690 18461
rect 20664 18429 20690 18432
rect 20664 18390 20690 18393
rect 20664 18361 20690 18364
rect 20526 18186 20552 18189
rect 20526 18157 20552 18160
rect 20388 15568 20414 15571
rect 20388 15539 20414 15542
rect 20256 11033 20362 11047
rect 20256 9383 20270 11033
rect 20342 10842 20368 10845
rect 20342 10813 20368 10816
rect 20296 10774 20322 10777
rect 20296 10745 20322 10748
rect 20302 10573 20316 10745
rect 20296 10570 20322 10573
rect 20296 10541 20322 10544
rect 20348 10539 20362 10813
rect 20342 10536 20368 10539
rect 20342 10507 20368 10510
rect 20250 9380 20276 9383
rect 20250 9351 20276 9354
rect 20394 8839 20408 15539
rect 20433 12628 20461 12632
rect 20433 12595 20434 12600
rect 20460 12595 20461 12600
rect 20480 12610 20506 12613
rect 20434 12581 20460 12584
rect 20480 12581 20506 12584
rect 20486 11865 20500 12581
rect 20480 11862 20506 11865
rect 20480 11833 20506 11836
rect 20434 10774 20460 10777
rect 20434 10745 20460 10748
rect 20440 9504 20454 10745
rect 20433 9500 20461 9504
rect 20461 9479 20500 9493
rect 20433 9467 20461 9472
rect 20434 9346 20460 9349
rect 20434 9317 20460 9320
rect 20250 8836 20276 8839
rect 20250 8807 20276 8810
rect 20388 8836 20414 8839
rect 20388 8807 20414 8810
rect 20204 8224 20230 8227
rect 20204 8195 20230 8198
rect 20210 8091 20224 8195
rect 20204 8088 20230 8091
rect 20204 8059 20230 8062
rect 20204 7816 20230 7819
rect 20204 7787 20230 7790
rect 20158 7000 20184 7003
rect 20158 6971 20184 6974
rect 19974 6932 20000 6935
rect 19974 6903 20000 6906
rect 19980 6119 19994 6903
rect 20210 6425 20224 7787
rect 20256 6697 20270 8807
rect 20342 8360 20368 8363
rect 20342 8331 20368 8334
rect 20348 8057 20362 8331
rect 20388 8326 20414 8329
rect 20388 8297 20414 8300
rect 20342 8054 20368 8057
rect 20342 8025 20368 8028
rect 20342 7510 20368 7513
rect 20342 7481 20368 7484
rect 20348 7173 20362 7481
rect 20342 7170 20368 7173
rect 20342 7141 20368 7144
rect 20348 6969 20362 7141
rect 20342 6966 20368 6969
rect 20342 6937 20368 6940
rect 20250 6694 20276 6697
rect 20250 6665 20276 6668
rect 20112 6422 20138 6425
rect 20112 6393 20138 6396
rect 20204 6422 20230 6425
rect 20204 6393 20230 6396
rect 20118 6217 20132 6393
rect 20118 6203 20178 6217
rect 20164 6119 20178 6203
rect 19882 6116 19908 6119
rect 19882 6087 19908 6090
rect 19974 6116 20000 6119
rect 19974 6087 20000 6090
rect 20158 6116 20184 6119
rect 20158 6087 20184 6090
rect 19330 5878 19356 5881
rect 19330 5849 19356 5852
rect 19836 5878 19862 5881
rect 19836 5849 19862 5852
rect 19842 5677 19856 5849
rect 19836 5674 19862 5677
rect 19836 5645 19862 5648
rect 19888 5575 19902 6087
rect 19980 5609 19994 6087
rect 20112 5844 20138 5847
rect 20112 5815 20138 5818
rect 19974 5606 20000 5609
rect 19974 5577 20000 5580
rect 19606 5572 19632 5575
rect 19606 5543 19632 5546
rect 19882 5572 19908 5575
rect 19882 5543 19908 5546
rect 19612 5031 19626 5543
rect 19888 5031 19902 5543
rect 20118 5371 20132 5815
rect 20112 5368 20138 5371
rect 20112 5339 20138 5342
rect 20164 5337 20178 6087
rect 20158 5334 20184 5337
rect 20158 5305 20184 5308
rect 19606 5028 19632 5031
rect 19606 4999 19632 5002
rect 19882 5028 19908 5031
rect 19882 4999 19908 5002
rect 19612 4827 19626 4999
rect 19606 4824 19632 4827
rect 19606 4795 19632 4798
rect 19612 4589 19626 4795
rect 19888 4793 19902 4999
rect 19882 4790 19908 4793
rect 19882 4761 19908 4764
rect 19606 4586 19632 4589
rect 19606 4557 19632 4560
rect 18640 3974 18666 3977
rect 18640 3945 18666 3948
rect 19192 3974 19218 3977
rect 19192 3945 19218 3948
rect 18646 1387 18660 3945
rect 20394 3943 20408 8297
rect 20440 8091 20454 9317
rect 20486 9043 20500 9479
rect 20532 9425 20546 18157
rect 20670 18087 20684 18361
rect 20664 18084 20690 18087
rect 20664 18055 20690 18058
rect 20670 17849 20684 18055
rect 20664 17846 20690 17849
rect 20664 17817 20690 17820
rect 20572 17200 20598 17203
rect 20572 17171 20598 17174
rect 20578 16999 20592 17171
rect 20572 16996 20598 16999
rect 20572 16967 20598 16970
rect 20578 16659 20592 16967
rect 20572 16656 20598 16659
rect 20572 16627 20598 16630
rect 20578 16183 20592 16627
rect 20572 16180 20598 16183
rect 20572 16151 20598 16154
rect 20578 15129 20592 16151
rect 20572 15126 20598 15129
rect 20572 15097 20598 15100
rect 20618 14106 20644 14109
rect 20618 14077 20644 14080
rect 20624 13939 20638 14077
rect 20618 13936 20644 13939
rect 20618 13907 20644 13910
rect 20716 11355 20730 18905
rect 20802 17302 20828 17305
rect 20802 17273 20828 17276
rect 20756 16758 20782 16761
rect 20756 16729 20782 16732
rect 20762 16115 20776 16729
rect 20808 16557 20822 17273
rect 20802 16554 20828 16557
rect 20802 16525 20828 16528
rect 20808 16251 20822 16525
rect 20802 16248 20828 16251
rect 20802 16219 20828 16222
rect 20756 16112 20782 16115
rect 20756 16083 20782 16086
rect 20762 15163 20776 16083
rect 20802 15670 20828 15673
rect 20802 15641 20828 15644
rect 20756 15160 20782 15163
rect 20756 15131 20782 15134
rect 20762 11865 20776 15131
rect 20808 15129 20822 15641
rect 20802 15126 20828 15129
rect 20802 15097 20828 15100
rect 20802 14004 20828 14007
rect 20802 13975 20828 13978
rect 20808 12987 20822 13975
rect 20854 13225 20868 22883
rect 21078 22436 21104 22439
rect 21078 22407 21104 22410
rect 21084 22201 21098 22407
rect 21078 22198 21104 22201
rect 21078 22169 21104 22172
rect 21084 21929 21098 22169
rect 21078 21926 21104 21929
rect 21078 21897 21104 21900
rect 21124 21892 21150 21895
rect 21124 21863 21150 21866
rect 20940 21110 20966 21113
rect 20940 21081 20966 21084
rect 20894 20260 20920 20263
rect 20894 20231 20920 20234
rect 20900 19957 20914 20231
rect 20946 20025 20960 21081
rect 21078 20804 21104 20807
rect 21078 20775 21104 20778
rect 21084 20535 21098 20775
rect 21130 20603 21144 21863
rect 21124 20600 21150 20603
rect 21124 20571 21150 20574
rect 21078 20532 21104 20535
rect 21078 20503 21104 20506
rect 20940 20022 20966 20025
rect 20940 19993 20966 19996
rect 20894 19954 20920 19957
rect 20894 19925 20920 19928
rect 20848 13222 20874 13225
rect 20848 13193 20874 13196
rect 20854 12987 20868 13193
rect 20802 12984 20828 12987
rect 20802 12955 20828 12958
rect 20848 12984 20874 12987
rect 20848 12955 20874 12958
rect 20854 12647 20868 12955
rect 20848 12644 20874 12647
rect 20848 12615 20874 12618
rect 20756 11862 20782 11865
rect 20756 11833 20782 11836
rect 20848 11862 20874 11865
rect 20848 11833 20874 11836
rect 20710 11352 20736 11355
rect 20710 11323 20736 11326
rect 20716 11047 20730 11323
rect 20716 11033 20776 11047
rect 20618 10672 20644 10675
rect 20618 10643 20644 10646
rect 20624 9757 20638 10643
rect 20618 9754 20644 9757
rect 20618 9725 20644 9728
rect 20572 9686 20598 9689
rect 20572 9657 20598 9660
rect 20578 9485 20592 9657
rect 20572 9482 20598 9485
rect 20572 9453 20598 9456
rect 20532 9411 20592 9425
rect 20526 9346 20552 9349
rect 20526 9317 20552 9320
rect 20532 9213 20546 9317
rect 20526 9210 20552 9213
rect 20526 9181 20552 9184
rect 20578 9145 20592 9411
rect 20664 9380 20690 9383
rect 20690 9354 20730 9357
rect 20664 9351 20730 9354
rect 20670 9343 20730 9351
rect 20572 9142 20598 9145
rect 20572 9113 20598 9116
rect 20480 9040 20506 9043
rect 20480 9011 20506 9014
rect 20716 8941 20730 9343
rect 20710 8938 20736 8941
rect 20710 8909 20736 8912
rect 20762 8133 20776 11033
rect 20716 8119 20776 8133
rect 20434 8088 20460 8091
rect 20434 8059 20460 8062
rect 20716 7411 20730 8119
rect 20756 8054 20782 8057
rect 20756 8025 20782 8028
rect 20762 7955 20776 8025
rect 20756 7952 20782 7955
rect 20756 7923 20782 7926
rect 20762 7547 20776 7923
rect 20756 7544 20782 7547
rect 20756 7515 20782 7518
rect 20710 7408 20736 7411
rect 20710 7379 20736 7382
rect 20571 6848 20599 6852
rect 20571 6815 20599 6820
rect 20578 6459 20592 6815
rect 20572 6456 20598 6459
rect 20572 6427 20598 6430
rect 20716 5915 20730 7379
rect 20710 5912 20736 5915
rect 20710 5883 20736 5886
rect 20854 5371 20868 11833
rect 20900 10811 20914 19925
rect 21084 19719 21098 20503
rect 21078 19716 21104 19719
rect 21078 19687 21104 19690
rect 21032 19478 21058 19481
rect 21032 19449 21058 19452
rect 21038 19141 21052 19449
rect 21084 19447 21098 19687
rect 21078 19444 21104 19447
rect 21078 19415 21104 19418
rect 21032 19138 21058 19141
rect 21032 19109 21058 19112
rect 20940 18594 20966 18597
rect 20940 18565 20966 18568
rect 20946 18412 20960 18565
rect 20939 18408 20967 18412
rect 20939 18375 20967 18380
rect 20946 15367 20960 18375
rect 21038 16217 21052 19109
rect 21078 18288 21104 18291
rect 21078 18259 21104 18262
rect 21084 18087 21098 18259
rect 21124 18186 21150 18189
rect 21124 18157 21150 18160
rect 21078 18084 21104 18087
rect 21078 18055 21104 18058
rect 21084 17815 21098 18055
rect 21078 17812 21104 17815
rect 21078 17783 21104 17786
rect 21084 17577 21098 17783
rect 21078 17574 21104 17577
rect 21078 17545 21104 17548
rect 21032 16214 21058 16217
rect 21032 16185 21058 16188
rect 20986 15840 21012 15843
rect 20986 15811 21012 15814
rect 20992 15760 21006 15811
rect 20985 15756 21013 15760
rect 20985 15723 21013 15728
rect 20992 15545 21006 15723
rect 21038 15639 21052 16185
rect 21032 15636 21058 15639
rect 21032 15607 21058 15610
rect 20992 15531 21052 15545
rect 20940 15364 20966 15367
rect 20940 15335 20966 15338
rect 21038 12987 21052 15531
rect 21130 14279 21144 18157
rect 21124 14276 21150 14279
rect 21124 14247 21150 14250
rect 21032 12984 21058 12987
rect 21032 12955 21058 12958
rect 21038 11047 21052 12955
rect 21176 11593 21190 24311
rect 21314 23799 21328 27099
rect 21544 26561 21558 33000
rect 21498 26553 21558 26561
rect 21492 26550 21558 26553
rect 21518 26547 21558 26550
rect 21492 26521 21518 26524
rect 21354 26006 21380 26009
rect 21354 25977 21380 25980
rect 21360 25635 21374 25977
rect 21544 25703 21558 26547
rect 22136 26448 22162 26451
rect 22136 26419 22162 26422
rect 22142 26043 22156 26419
rect 22136 26040 22162 26043
rect 22136 26011 22162 26014
rect 21584 25972 21610 25975
rect 21584 25943 21610 25946
rect 21538 25700 21564 25703
rect 21538 25671 21564 25674
rect 21354 25632 21380 25635
rect 21354 25603 21380 25606
rect 21446 25632 21472 25635
rect 21446 25603 21472 25606
rect 21308 23796 21334 23799
rect 21308 23767 21334 23770
rect 21216 23592 21242 23595
rect 21216 23563 21242 23566
rect 21222 23323 21236 23563
rect 21262 23490 21288 23493
rect 21262 23461 21288 23464
rect 21216 23320 21242 23323
rect 21216 23291 21242 23294
rect 21268 23085 21282 23461
rect 21262 23082 21288 23085
rect 21262 23053 21288 23056
rect 21314 23017 21328 23767
rect 21360 23527 21374 25603
rect 21400 24918 21426 24921
rect 21400 24889 21426 24892
rect 21406 24071 21420 24889
rect 21400 24068 21426 24071
rect 21400 24039 21426 24042
rect 21452 23833 21466 25603
rect 21544 24887 21558 25671
rect 21590 25635 21604 25943
rect 21584 25632 21610 25635
rect 21584 25603 21610 25606
rect 21676 25156 21702 25159
rect 21676 25127 21702 25130
rect 21538 24884 21564 24887
rect 21538 24855 21564 24858
rect 21682 24615 21696 25127
rect 21906 25122 21932 25125
rect 21906 25093 21932 25096
rect 21912 24649 21926 25093
rect 21906 24646 21932 24649
rect 21906 24617 21932 24620
rect 21676 24612 21702 24615
rect 21676 24583 21702 24586
rect 21682 24105 21696 24583
rect 21676 24102 21702 24105
rect 21676 24073 21702 24076
rect 21682 23909 21696 24073
rect 21912 24045 21926 24617
rect 21998 24578 22024 24581
rect 21998 24549 22024 24552
rect 22004 24521 22018 24549
rect 22004 24507 22110 24521
rect 22096 24377 22110 24507
rect 22832 24411 22846 33000
rect 22970 32968 23168 32982
rect 22872 25904 22898 25907
rect 22872 25875 22898 25878
rect 22878 25703 22892 25875
rect 22872 25700 22898 25703
rect 22872 25671 22898 25674
rect 22826 24408 22852 24411
rect 22826 24379 22852 24382
rect 22090 24374 22116 24377
rect 22090 24345 22116 24348
rect 21912 24037 21972 24045
rect 21912 24034 21978 24037
rect 21912 24031 21952 24034
rect 21952 24005 21978 24008
rect 21584 23898 21610 23901
rect 21682 23895 21742 23909
rect 21584 23869 21610 23872
rect 21446 23830 21472 23833
rect 21446 23801 21472 23804
rect 21492 23728 21518 23731
rect 21492 23699 21518 23702
rect 21400 23558 21426 23561
rect 21400 23529 21426 23532
rect 21354 23524 21380 23527
rect 21354 23495 21380 23498
rect 21406 23433 21420 23529
rect 21360 23419 21420 23433
rect 21360 23289 21374 23419
rect 21498 23323 21512 23699
rect 21590 23459 21604 23869
rect 21676 23864 21702 23867
rect 21676 23835 21702 23838
rect 21584 23456 21610 23459
rect 21584 23427 21610 23430
rect 21492 23320 21518 23323
rect 21492 23291 21518 23294
rect 21354 23286 21380 23289
rect 21354 23257 21380 23260
rect 21216 23014 21242 23017
rect 21216 22985 21242 22988
rect 21308 23014 21334 23017
rect 21308 22985 21334 22988
rect 21222 22915 21236 22985
rect 21216 22912 21242 22915
rect 21216 22883 21242 22886
rect 21360 22439 21374 23257
rect 21590 22983 21604 23427
rect 21682 23085 21696 23835
rect 21728 23561 21742 23895
rect 21958 23569 21972 24005
rect 21722 23558 21748 23561
rect 21958 23555 22064 23569
rect 21722 23529 21748 23532
rect 21952 23524 21978 23527
rect 21952 23495 21978 23498
rect 21676 23082 21702 23085
rect 21676 23053 21702 23056
rect 21584 22980 21610 22983
rect 21584 22951 21610 22954
rect 21630 22980 21656 22983
rect 21630 22951 21656 22954
rect 21538 22776 21564 22779
rect 21538 22747 21564 22750
rect 21354 22436 21380 22439
rect 21354 22407 21380 22410
rect 21544 22405 21558 22747
rect 21636 22439 21650 22951
rect 21958 22745 21972 23495
rect 22050 23493 22064 23555
rect 22044 23490 22070 23493
rect 22044 23461 22070 23464
rect 22044 23184 22070 23187
rect 22044 23155 22070 23158
rect 22050 22983 22064 23155
rect 22044 22980 22070 22983
rect 22044 22951 22070 22954
rect 21952 22742 21978 22745
rect 21952 22713 21978 22716
rect 22096 22711 22110 24345
rect 22688 23592 22714 23595
rect 22688 23563 22714 23566
rect 22694 23085 22708 23563
rect 22688 23082 22714 23085
rect 22688 23053 22714 23056
rect 22832 22983 22846 24379
rect 22970 24377 22984 32968
rect 23154 32953 23168 32968
rect 23200 32953 23214 33000
rect 23154 32939 23214 32953
rect 23010 26006 23036 26009
rect 23010 25977 23036 25980
rect 23286 26006 23312 26009
rect 23286 25977 23312 25980
rect 23332 26006 23358 26009
rect 23332 25977 23358 25980
rect 23016 25805 23030 25977
rect 23010 25802 23036 25805
rect 23010 25773 23036 25776
rect 23102 25700 23128 25703
rect 23102 25671 23128 25674
rect 23108 25397 23122 25671
rect 23292 25431 23306 25977
rect 23338 25465 23352 25977
rect 23378 25972 23404 25975
rect 23378 25943 23404 25946
rect 23332 25462 23358 25465
rect 23332 25433 23358 25436
rect 23286 25428 23312 25431
rect 23286 25399 23312 25402
rect 23102 25394 23128 25397
rect 23102 25365 23128 25368
rect 23108 25261 23122 25365
rect 23102 25258 23128 25261
rect 23102 25229 23128 25232
rect 22964 24374 22990 24377
rect 22964 24345 22990 24348
rect 23240 24374 23266 24377
rect 23240 24345 23266 24348
rect 22918 24340 22944 24343
rect 22918 24311 22944 24314
rect 22924 24173 22938 24311
rect 22918 24170 22944 24173
rect 22918 24141 22944 24144
rect 23246 24071 23260 24345
rect 23292 24309 23306 25399
rect 23338 24717 23352 25433
rect 23332 24714 23358 24717
rect 23332 24685 23358 24688
rect 23384 24377 23398 25943
rect 23654 25734 23680 25737
rect 23654 25705 23680 25708
rect 23660 25533 23674 25705
rect 23654 25530 23680 25533
rect 23654 25501 23680 25504
rect 23562 25360 23588 25363
rect 23562 25331 23588 25334
rect 23568 24445 23582 25331
rect 23660 24717 23674 25501
rect 23936 25159 23950 33000
rect 24028 32953 24042 33000
rect 24074 32968 24134 32982
rect 24074 32953 24088 32968
rect 24028 32939 24088 32953
rect 23930 25156 23956 25159
rect 23930 25127 23956 25130
rect 23654 24714 23680 24717
rect 23654 24685 23680 24688
rect 23936 24615 23950 25127
rect 23930 24612 23956 24615
rect 23930 24583 23956 24586
rect 24068 24578 24094 24581
rect 24068 24549 24094 24552
rect 23562 24442 23588 24445
rect 23562 24413 23588 24416
rect 23470 24408 23496 24411
rect 23430 24382 23470 24385
rect 23430 24379 23496 24382
rect 23378 24374 23404 24377
rect 23378 24345 23404 24348
rect 23430 24371 23490 24379
rect 24074 24377 24088 24549
rect 24120 24411 24134 32968
rect 24114 24408 24140 24411
rect 24114 24379 24140 24382
rect 23746 24374 23772 24377
rect 23286 24306 23312 24309
rect 23286 24277 23312 24280
rect 23240 24068 23266 24071
rect 23240 24039 23266 24042
rect 22826 22980 22852 22983
rect 22826 22951 22852 22954
rect 23194 22980 23220 22983
rect 23194 22951 23220 22954
rect 22090 22708 22116 22711
rect 22090 22679 22116 22682
rect 21630 22436 21656 22439
rect 21630 22407 21656 22410
rect 23056 22436 23082 22439
rect 23056 22407 23082 22410
rect 21538 22402 21564 22405
rect 21538 22373 21564 22376
rect 21307 22352 21335 22356
rect 21307 22319 21335 22324
rect 21314 22235 21328 22319
rect 21308 22232 21334 22235
rect 21268 22212 21308 22226
rect 21216 21382 21242 21385
rect 21216 21353 21242 21356
rect 21222 20739 21236 21353
rect 21216 20736 21242 20739
rect 21216 20707 21242 20710
rect 21222 20569 21236 20707
rect 21216 20566 21242 20569
rect 21216 20537 21242 20540
rect 21268 20509 21282 22212
rect 21308 22203 21334 22206
rect 21446 21858 21472 21861
rect 21446 21829 21472 21832
rect 21452 21725 21466 21829
rect 21446 21722 21472 21725
rect 21446 21693 21472 21696
rect 21446 20770 21472 20773
rect 21446 20741 21472 20744
rect 21354 20566 21380 20569
rect 21354 20537 21380 20540
rect 21222 20495 21282 20509
rect 21222 17747 21236 20495
rect 21262 19716 21288 19719
rect 21262 19687 21288 19690
rect 21268 19175 21282 19687
rect 21360 19685 21374 20537
rect 21452 20365 21466 20741
rect 21446 20362 21472 20365
rect 21446 20333 21472 20336
rect 21452 19821 21466 20333
rect 21446 19818 21472 19821
rect 21446 19789 21472 19792
rect 21354 19682 21380 19685
rect 21354 19653 21380 19656
rect 21308 19512 21334 19515
rect 21308 19483 21334 19486
rect 21262 19172 21288 19175
rect 21262 19143 21288 19146
rect 21262 18560 21288 18563
rect 21262 18531 21288 18534
rect 21216 17744 21242 17747
rect 21216 17715 21242 17718
rect 21216 17574 21242 17577
rect 21216 17545 21242 17548
rect 21222 17033 21236 17545
rect 21216 17030 21242 17033
rect 21216 17001 21242 17004
rect 21268 16829 21282 18531
rect 21314 18393 21328 19483
rect 21360 19481 21374 19653
rect 21354 19478 21380 19481
rect 21354 19449 21380 19452
rect 21354 19172 21380 19175
rect 21354 19143 21380 19146
rect 21360 18971 21374 19143
rect 21354 18968 21380 18971
rect 21354 18939 21380 18942
rect 21354 18560 21380 18563
rect 21354 18531 21380 18534
rect 21308 18390 21334 18393
rect 21308 18361 21334 18364
rect 21360 18189 21374 18531
rect 21354 18186 21380 18189
rect 21354 18157 21380 18160
rect 21446 18186 21472 18189
rect 21446 18157 21472 18160
rect 21452 18053 21466 18157
rect 21446 18050 21472 18053
rect 21446 18021 21472 18024
rect 21354 17880 21380 17883
rect 21354 17851 21380 17854
rect 21360 17747 21374 17851
rect 21354 17744 21380 17747
rect 21354 17715 21380 17718
rect 21262 16826 21288 16829
rect 21262 16797 21288 16800
rect 21308 16758 21334 16761
rect 21308 16729 21334 16732
rect 21261 16640 21289 16644
rect 21261 16607 21289 16612
rect 21216 13188 21242 13191
rect 21216 13159 21242 13162
rect 21222 12851 21236 13159
rect 21216 12848 21242 12851
rect 21216 12819 21242 12822
rect 21222 12681 21236 12819
rect 21216 12678 21242 12681
rect 21216 12649 21242 12652
rect 21170 11590 21196 11593
rect 21170 11561 21196 11564
rect 21222 11261 21236 12649
rect 21176 11247 21236 11261
rect 21176 11219 21190 11247
rect 21170 11216 21196 11219
rect 21170 11187 21196 11190
rect 21176 11049 21190 11187
rect 20946 11033 21052 11047
rect 21170 11046 21196 11049
rect 20894 10808 20920 10811
rect 20894 10779 20920 10782
rect 20900 8295 20914 10779
rect 20946 9232 20960 11033
rect 21170 11017 21196 11020
rect 21176 10675 21190 11017
rect 21216 10978 21242 10981
rect 21216 10949 21242 10952
rect 21222 10777 21236 10949
rect 21216 10774 21242 10777
rect 21216 10745 21242 10748
rect 21170 10672 21196 10675
rect 21170 10643 21196 10646
rect 20939 9228 20967 9232
rect 20939 9195 20967 9200
rect 20894 8292 20920 8295
rect 20894 8263 20920 8266
rect 20946 7785 20960 9195
rect 21268 8677 21282 16607
rect 21314 16455 21328 16729
rect 21360 16644 21374 17715
rect 21452 17245 21466 18021
rect 21492 17846 21518 17849
rect 21492 17817 21518 17820
rect 21406 17231 21466 17245
rect 21406 16701 21420 17231
rect 21446 17200 21472 17203
rect 21446 17171 21472 17174
rect 21452 16761 21466 17171
rect 21498 16999 21512 17817
rect 21544 16999 21558 22373
rect 21636 22201 21650 22407
rect 22734 22368 22760 22371
rect 22734 22339 22760 22342
rect 23010 22368 23036 22371
rect 23010 22339 23036 22342
rect 21630 22198 21656 22201
rect 21630 22169 21656 22172
rect 21636 21895 21650 22169
rect 22642 22096 22668 22099
rect 22642 22067 22668 22070
rect 22648 21895 22662 22067
rect 22740 21929 22754 22339
rect 23016 22235 23030 22339
rect 23010 22232 23036 22235
rect 23010 22203 23036 22206
rect 23062 21997 23076 22407
rect 23056 21994 23082 21997
rect 23056 21965 23082 21968
rect 22734 21926 22760 21929
rect 22734 21897 22760 21900
rect 21630 21892 21656 21895
rect 21630 21863 21656 21866
rect 22504 21892 22530 21895
rect 22642 21892 22668 21895
rect 22530 21872 22570 21886
rect 22504 21863 22530 21866
rect 21636 21385 21650 21863
rect 22320 21858 22346 21861
rect 22320 21829 22346 21832
rect 21676 21722 21702 21725
rect 21676 21693 21702 21696
rect 21630 21382 21656 21385
rect 21630 21353 21656 21356
rect 21584 19716 21610 19719
rect 21584 19687 21610 19690
rect 21590 18189 21604 19687
rect 21629 18612 21657 18616
rect 21629 18579 21657 18584
rect 21636 18393 21650 18579
rect 21630 18390 21656 18393
rect 21630 18361 21656 18364
rect 21584 18186 21610 18189
rect 21584 18157 21610 18160
rect 21636 18129 21650 18361
rect 21590 18115 21650 18129
rect 21492 16996 21518 16999
rect 21492 16967 21518 16970
rect 21538 16996 21564 16999
rect 21538 16967 21564 16970
rect 21446 16758 21472 16761
rect 21446 16729 21472 16732
rect 21406 16687 21512 16701
rect 21353 16640 21381 16644
rect 21353 16607 21381 16612
rect 21308 16452 21334 16455
rect 21308 16423 21334 16426
rect 21314 15630 21328 16423
rect 21400 15636 21426 15639
rect 21314 15616 21400 15630
rect 21400 15607 21426 15610
rect 21354 14310 21380 14313
rect 21354 14281 21380 14284
rect 21360 14109 21374 14281
rect 21354 14106 21380 14109
rect 21354 14077 21380 14080
rect 21360 13429 21374 14077
rect 21406 14049 21420 15607
rect 21498 14389 21512 16687
rect 21544 14823 21558 16967
rect 21538 14820 21564 14823
rect 21538 14791 21564 14794
rect 21498 14375 21558 14389
rect 21492 14344 21518 14347
rect 21492 14315 21518 14318
rect 21446 14208 21472 14211
rect 21446 14179 21472 14182
rect 21452 14109 21466 14179
rect 21446 14106 21472 14109
rect 21446 14077 21472 14080
rect 21498 14075 21512 14315
rect 21492 14072 21518 14075
rect 21406 14035 21466 14049
rect 21492 14043 21518 14046
rect 21400 13460 21426 13463
rect 21400 13431 21426 13434
rect 21354 13426 21380 13429
rect 21354 13397 21380 13400
rect 21406 10989 21420 13431
rect 21452 11899 21466 14035
rect 21492 14004 21518 14007
rect 21492 13975 21518 13978
rect 21498 13701 21512 13975
rect 21492 13698 21518 13701
rect 21492 13669 21518 13672
rect 21498 12307 21512 13669
rect 21544 13191 21558 14375
rect 21590 13463 21604 18115
rect 21630 18084 21656 18087
rect 21682 18078 21696 21693
rect 22326 18631 22340 21829
rect 22504 21824 22530 21827
rect 22504 21795 22530 21798
rect 22458 21722 22484 21725
rect 22458 21693 22484 21696
rect 22366 18662 22392 18665
rect 22366 18633 22392 18636
rect 21952 18628 21978 18631
rect 21952 18599 21978 18602
rect 22090 18628 22116 18631
rect 22090 18599 22116 18602
rect 22320 18628 22346 18631
rect 22320 18599 22346 18602
rect 21958 18461 21972 18599
rect 21952 18458 21978 18461
rect 21952 18429 21978 18432
rect 22096 18189 22110 18599
rect 22090 18186 22116 18189
rect 22090 18157 22116 18160
rect 22326 18155 22340 18599
rect 22320 18152 22346 18155
rect 22320 18123 22346 18126
rect 21656 18064 21696 18078
rect 21630 18055 21656 18058
rect 22372 17917 22386 18633
rect 22464 18548 22478 21693
rect 22510 20841 22524 21795
rect 22556 21725 22570 21872
rect 22642 21863 22668 21866
rect 23010 21892 23036 21895
rect 23010 21863 23036 21866
rect 22550 21722 22576 21725
rect 22550 21693 22576 21696
rect 22642 21008 22668 21011
rect 22642 20979 22668 20982
rect 22504 20838 22530 20841
rect 22504 20809 22530 20812
rect 22648 20807 22662 20979
rect 22642 20804 22668 20807
rect 22642 20775 22668 20778
rect 22688 20770 22714 20773
rect 22688 20741 22714 20744
rect 22872 20770 22898 20773
rect 22872 20741 22898 20744
rect 22550 20736 22576 20739
rect 22550 20707 22576 20710
rect 22596 20736 22622 20739
rect 22596 20707 22622 20710
rect 22556 20603 22570 20707
rect 22550 20600 22576 20603
rect 22550 20571 22576 20574
rect 22602 19549 22616 20707
rect 22642 20566 22668 20569
rect 22642 20537 22668 20540
rect 22648 20263 22662 20537
rect 22694 20501 22708 20741
rect 22688 20498 22714 20501
rect 22688 20469 22714 20472
rect 22642 20260 22668 20263
rect 22642 20231 22668 20234
rect 22596 19546 22622 19549
rect 22596 19517 22622 19520
rect 22596 19478 22622 19481
rect 22596 19449 22622 19452
rect 22602 18733 22616 19449
rect 22648 19379 22662 20231
rect 22688 20022 22714 20025
rect 22688 19993 22714 19996
rect 22694 19787 22708 19993
rect 22688 19784 22714 19787
rect 22688 19755 22714 19758
rect 22694 19421 22708 19755
rect 22734 19648 22760 19651
rect 22734 19619 22760 19622
rect 22740 19481 22754 19619
rect 22780 19546 22806 19549
rect 22780 19517 22806 19520
rect 22734 19478 22760 19481
rect 22734 19449 22760 19452
rect 22694 19407 22754 19421
rect 22642 19376 22668 19379
rect 22642 19347 22668 19350
rect 22596 18730 22622 18733
rect 22596 18701 22622 18704
rect 22457 18544 22485 18548
rect 22457 18511 22485 18516
rect 22366 17914 22392 17917
rect 22366 17885 22392 17888
rect 22458 17744 22484 17747
rect 22458 17715 22484 17718
rect 22464 17577 22478 17715
rect 22458 17574 22484 17577
rect 22458 17545 22484 17548
rect 22043 17524 22071 17528
rect 21630 17506 21656 17509
rect 22043 17491 22044 17496
rect 21630 17477 21656 17480
rect 22070 17491 22071 17496
rect 22688 17506 22714 17509
rect 22044 17477 22070 17480
rect 22688 17477 22714 17480
rect 21636 15673 21650 17477
rect 22694 16965 22708 17477
rect 22688 16962 22714 16965
rect 22688 16933 22714 16936
rect 21676 16928 21702 16931
rect 22694 16916 22708 16933
rect 21676 16899 21702 16902
rect 22687 16912 22715 16916
rect 21682 16795 21696 16899
rect 22687 16879 22715 16884
rect 22688 16826 22714 16829
rect 22688 16797 22714 16800
rect 21676 16792 21702 16795
rect 21676 16763 21702 16766
rect 22694 16761 22708 16797
rect 22688 16758 22714 16761
rect 22688 16729 22714 16732
rect 21906 16690 21932 16693
rect 21906 16661 21932 16664
rect 21860 16112 21886 16115
rect 21860 16083 21886 16086
rect 21866 15741 21880 16083
rect 21860 15738 21886 15741
rect 21860 15709 21886 15712
rect 21912 15673 21926 16661
rect 21630 15670 21656 15673
rect 21630 15641 21656 15644
rect 21722 15670 21748 15673
rect 21722 15641 21748 15644
rect 21906 15670 21932 15673
rect 21906 15641 21932 15644
rect 21728 15197 21742 15641
rect 21722 15194 21748 15197
rect 21722 15165 21748 15168
rect 21584 13460 21610 13463
rect 21584 13431 21610 13434
rect 21912 13191 21926 15641
rect 22642 15466 22668 15469
rect 22642 15437 22668 15440
rect 22044 14820 22070 14823
rect 22044 14791 22070 14794
rect 21538 13188 21564 13191
rect 21538 13159 21564 13162
rect 21906 13188 21932 13191
rect 21906 13159 21932 13162
rect 21492 12304 21518 12307
rect 21492 12275 21518 12278
rect 21446 11896 21472 11899
rect 21446 11867 21472 11870
rect 21406 10981 21466 10989
rect 21406 10978 21472 10981
rect 21406 10975 21446 10978
rect 21353 10860 21381 10864
rect 21353 10827 21381 10832
rect 21360 10811 21374 10827
rect 21354 10808 21380 10811
rect 21354 10779 21380 10782
rect 21406 9451 21420 10975
rect 21446 10949 21472 10952
rect 21400 9448 21426 9451
rect 21400 9419 21426 9422
rect 21354 9414 21380 9417
rect 21354 9385 21380 9388
rect 21360 9300 21374 9385
rect 21353 9296 21381 9300
rect 21353 9263 21381 9268
rect 21222 8663 21282 8677
rect 21032 8122 21058 8125
rect 21032 8093 21058 8096
rect 20986 7986 21012 7989
rect 20986 7957 21012 7960
rect 20940 7782 20966 7785
rect 20940 7753 20966 7756
rect 20992 7513 21006 7957
rect 21038 7547 21052 8093
rect 21078 8054 21104 8057
rect 21078 8025 21104 8028
rect 21084 7717 21098 8025
rect 21078 7714 21104 7717
rect 21078 7685 21104 7688
rect 21084 7547 21098 7685
rect 21032 7544 21058 7547
rect 21032 7515 21058 7518
rect 21078 7544 21104 7547
rect 21078 7515 21104 7518
rect 20986 7510 21012 7513
rect 20986 7481 21012 7484
rect 21078 7306 21104 7309
rect 21078 7277 21104 7280
rect 21084 6969 21098 7277
rect 21222 7139 21236 8663
rect 21262 8598 21288 8601
rect 21262 8569 21288 8572
rect 21308 8598 21334 8601
rect 21308 8569 21334 8572
rect 21268 8363 21282 8569
rect 21262 8360 21288 8363
rect 21262 8331 21288 8334
rect 21314 8295 21328 8569
rect 21308 8292 21334 8295
rect 21308 8263 21334 8266
rect 21314 8125 21328 8263
rect 21360 8125 21374 9263
rect 21308 8122 21334 8125
rect 21308 8093 21334 8096
rect 21354 8122 21380 8125
rect 21354 8093 21380 8096
rect 21406 7445 21420 9419
rect 21544 8635 21558 13159
rect 21629 12696 21657 12700
rect 21629 12663 21657 12668
rect 21636 12647 21650 12663
rect 21630 12644 21656 12647
rect 21630 12615 21656 12618
rect 21584 12066 21610 12069
rect 21584 12037 21610 12040
rect 21590 11831 21604 12037
rect 21630 11862 21656 11865
rect 21630 11833 21656 11836
rect 21676 11862 21702 11865
rect 21676 11833 21702 11836
rect 21722 11862 21748 11865
rect 21722 11833 21748 11836
rect 21584 11828 21610 11831
rect 21584 11799 21610 11802
rect 21636 11047 21650 11833
rect 21682 11389 21696 11833
rect 21728 11763 21742 11833
rect 21722 11760 21748 11763
rect 21722 11731 21748 11734
rect 21676 11386 21702 11389
rect 21676 11357 21702 11360
rect 21636 11033 21696 11047
rect 21538 8632 21564 8635
rect 21538 8603 21564 8606
rect 21544 7785 21558 8603
rect 21630 8598 21656 8601
rect 21630 8569 21656 8572
rect 21636 8057 21650 8569
rect 21630 8054 21656 8057
rect 21630 8025 21656 8028
rect 21636 7785 21650 8025
rect 21538 7782 21564 7785
rect 21538 7753 21564 7756
rect 21630 7782 21656 7785
rect 21630 7753 21656 7756
rect 21446 7748 21472 7751
rect 21446 7719 21472 7722
rect 21452 7581 21466 7719
rect 21682 7683 21696 11033
rect 21728 9621 21742 11731
rect 21722 9618 21748 9621
rect 21722 9589 21748 9592
rect 21998 9346 22024 9349
rect 21998 9317 22024 9320
rect 21952 9312 21978 9315
rect 21952 9283 21978 9286
rect 21676 7680 21702 7683
rect 21676 7651 21702 7654
rect 21446 7578 21472 7581
rect 21446 7549 21472 7552
rect 21400 7442 21426 7445
rect 21400 7413 21426 7416
rect 21400 7272 21426 7275
rect 21400 7243 21426 7246
rect 21308 7170 21334 7173
rect 21308 7141 21334 7144
rect 21124 7136 21150 7139
rect 21124 7107 21150 7110
rect 21216 7136 21242 7139
rect 21216 7107 21242 7110
rect 21130 7037 21144 7107
rect 21124 7034 21150 7037
rect 21124 7005 21150 7008
rect 21314 7003 21328 7141
rect 21308 7000 21334 7003
rect 21308 6971 21334 6974
rect 21078 6966 21104 6969
rect 21078 6937 21104 6940
rect 21354 6966 21380 6969
rect 21354 6937 21380 6940
rect 21084 6663 21098 6937
rect 21261 6712 21289 6716
rect 21261 6679 21289 6684
rect 21268 6663 21282 6679
rect 21360 6663 21374 6937
rect 21078 6660 21104 6663
rect 21078 6631 21104 6634
rect 21262 6660 21288 6663
rect 21262 6631 21288 6634
rect 21354 6660 21380 6663
rect 21354 6631 21380 6634
rect 21084 6425 21098 6631
rect 21124 6626 21150 6629
rect 21124 6597 21150 6600
rect 21078 6422 21104 6425
rect 21078 6393 21104 6396
rect 20848 5368 20874 5371
rect 20848 5339 20874 5342
rect 20854 5235 20868 5339
rect 21084 5337 21098 6393
rect 21078 5334 21104 5337
rect 21078 5305 21104 5308
rect 20848 5232 20874 5235
rect 20848 5203 20874 5206
rect 21084 5065 21098 5305
rect 21078 5062 21104 5065
rect 21078 5033 21104 5036
rect 21084 4793 21098 5033
rect 21130 4827 21144 6597
rect 21268 5821 21282 6631
rect 21307 6508 21335 6512
rect 21307 6475 21335 6480
rect 21314 6459 21328 6475
rect 21308 6456 21334 6459
rect 21308 6427 21334 6430
rect 21314 6153 21328 6427
rect 21360 6425 21374 6631
rect 21354 6422 21380 6425
rect 21354 6393 21380 6396
rect 21308 6150 21334 6153
rect 21308 6121 21334 6124
rect 21268 5807 21328 5821
rect 21314 5371 21328 5807
rect 21308 5368 21334 5371
rect 21308 5339 21334 5342
rect 21360 5337 21374 6393
rect 21406 6217 21420 7243
rect 21446 7136 21472 7139
rect 21446 7107 21472 7110
rect 21452 6629 21466 7107
rect 21958 6988 21972 9283
rect 22004 9145 22018 9317
rect 21998 9142 22024 9145
rect 21998 9113 22024 9116
rect 22004 8805 22018 9113
rect 22050 8907 22064 14791
rect 22320 13834 22346 13837
rect 22320 13805 22346 13808
rect 22274 12916 22300 12919
rect 22274 12887 22300 12890
rect 22280 12749 22294 12887
rect 22274 12746 22300 12749
rect 22274 12717 22300 12720
rect 22090 12100 22116 12103
rect 22090 12071 22116 12074
rect 22096 11049 22110 12071
rect 22090 11046 22116 11049
rect 22090 11017 22116 11020
rect 22326 9893 22340 13805
rect 22648 12953 22662 15437
rect 22694 14381 22708 16729
rect 22688 14378 22714 14381
rect 22688 14349 22714 14352
rect 22694 13837 22708 14349
rect 22688 13834 22714 13837
rect 22688 13805 22714 13808
rect 22642 12950 22668 12953
rect 22642 12921 22668 12924
rect 22596 12848 22622 12851
rect 22596 12819 22622 12822
rect 22412 12678 22438 12681
rect 22412 12649 22438 12652
rect 22320 9890 22346 9893
rect 22320 9861 22346 9864
rect 22182 9856 22208 9859
rect 22182 9827 22208 9830
rect 22090 9652 22116 9655
rect 22090 9623 22116 9626
rect 22044 8904 22070 8907
rect 22044 8875 22070 8878
rect 21998 8802 22024 8805
rect 21998 8773 22024 8776
rect 22004 8295 22018 8773
rect 21998 8292 22024 8295
rect 21998 8263 22024 8266
rect 21951 6984 21979 6988
rect 21951 6951 21979 6956
rect 21446 6626 21472 6629
rect 21446 6597 21472 6600
rect 21452 6580 21466 6597
rect 21445 6576 21473 6580
rect 21445 6543 21473 6548
rect 21406 6203 21466 6217
rect 21354 5334 21380 5337
rect 21354 5305 21380 5308
rect 21360 5031 21374 5305
rect 21354 5028 21380 5031
rect 21452 5016 21466 6203
rect 21958 5541 21972 6951
rect 22096 6901 22110 9623
rect 22188 9417 22202 9827
rect 22320 9720 22346 9723
rect 22320 9691 22346 9694
rect 22182 9414 22208 9417
rect 22182 9385 22208 9388
rect 22182 8836 22208 8839
rect 22182 8807 22208 8810
rect 22188 8601 22202 8807
rect 22182 8598 22208 8601
rect 22182 8569 22208 8572
rect 22228 8598 22254 8601
rect 22228 8569 22254 8572
rect 22136 8530 22162 8533
rect 22136 8501 22162 8504
rect 22142 8023 22156 8501
rect 22136 8020 22162 8023
rect 22136 7991 22162 7994
rect 22136 7952 22162 7955
rect 22136 7923 22162 7926
rect 22142 7751 22156 7923
rect 22188 7751 22202 8569
rect 22234 8295 22248 8569
rect 22228 8292 22254 8295
rect 22228 8263 22254 8266
rect 22234 7955 22248 8263
rect 22274 8020 22300 8023
rect 22274 7991 22300 7994
rect 22228 7952 22254 7955
rect 22228 7923 22254 7926
rect 22280 7819 22294 7991
rect 22274 7816 22300 7819
rect 22274 7787 22300 7790
rect 22136 7748 22162 7751
rect 22136 7719 22162 7722
rect 22182 7748 22208 7751
rect 22182 7719 22208 7722
rect 22142 7207 22156 7719
rect 22188 7241 22202 7719
rect 22182 7238 22208 7241
rect 22182 7209 22208 7212
rect 22136 7204 22162 7207
rect 22136 7175 22162 7178
rect 22090 6898 22116 6901
rect 22090 6869 22116 6872
rect 22280 5643 22294 7787
rect 22274 5640 22300 5643
rect 22274 5611 22300 5614
rect 22136 5572 22162 5575
rect 22136 5543 22162 5546
rect 22274 5572 22300 5575
rect 22274 5543 22300 5546
rect 21952 5538 21978 5541
rect 21952 5509 21978 5512
rect 22142 5133 22156 5543
rect 22280 5405 22294 5543
rect 22326 5507 22340 9691
rect 22418 9368 22432 12649
rect 22602 12137 22616 12819
rect 22648 12681 22662 12921
rect 22642 12678 22668 12681
rect 22642 12649 22668 12652
rect 22596 12134 22622 12137
rect 22596 12105 22622 12108
rect 22740 11047 22754 19407
rect 22786 19277 22800 19517
rect 22826 19376 22852 19379
rect 22826 19347 22852 19350
rect 22780 19274 22806 19277
rect 22780 19245 22806 19248
rect 22832 18699 22846 19347
rect 22826 18696 22852 18699
rect 22826 18667 22852 18670
rect 22780 18390 22806 18393
rect 22780 18361 22806 18364
rect 22786 17849 22800 18361
rect 22780 17846 22806 17849
rect 22780 17817 22806 17820
rect 22786 17543 22800 17817
rect 22780 17540 22806 17543
rect 22780 17511 22806 17514
rect 22780 16758 22806 16761
rect 22780 16729 22806 16732
rect 22786 16217 22800 16729
rect 22780 16214 22806 16217
rect 22780 16185 22806 16188
rect 22832 16157 22846 18667
rect 22786 16143 22846 16157
rect 22786 13021 22800 16143
rect 22826 15568 22852 15571
rect 22826 15539 22852 15542
rect 22832 15401 22846 15539
rect 22826 15398 22852 15401
rect 22826 15369 22852 15372
rect 22878 15367 22892 20741
rect 22918 20566 22944 20569
rect 22918 20537 22944 20540
rect 22924 19976 22938 20537
rect 22917 19972 22945 19976
rect 22917 19939 22945 19944
rect 22964 19954 22990 19957
rect 22924 19568 22938 19939
rect 22964 19925 22990 19928
rect 22970 19651 22984 19925
rect 22964 19648 22990 19651
rect 22964 19619 22990 19622
rect 22917 19564 22945 19568
rect 22917 19531 22945 19536
rect 22970 19515 22984 19619
rect 22964 19512 22990 19515
rect 22964 19483 22990 19486
rect 22918 19478 22944 19481
rect 22918 19449 22944 19452
rect 22924 18835 22938 19449
rect 22964 19444 22990 19447
rect 22964 19415 22990 19418
rect 22970 18971 22984 19415
rect 22964 18968 22990 18971
rect 22964 18939 22990 18942
rect 22918 18832 22944 18835
rect 22918 18803 22944 18806
rect 22924 17645 22938 18803
rect 22970 18359 22984 18939
rect 22964 18356 22990 18359
rect 22964 18327 22990 18330
rect 22964 17880 22990 17883
rect 22964 17851 22990 17854
rect 22918 17642 22944 17645
rect 22918 17613 22944 17616
rect 22918 16792 22944 16795
rect 22918 16763 22944 16766
rect 22924 16557 22938 16763
rect 22918 16554 22944 16557
rect 22918 16525 22944 16528
rect 22970 15843 22984 17851
rect 23016 16829 23030 21863
rect 23200 21861 23214 22951
rect 23246 21895 23260 24039
rect 23430 23569 23444 24371
rect 23746 24345 23772 24348
rect 24068 24374 24094 24377
rect 24068 24345 24094 24348
rect 23608 24000 23634 24003
rect 23608 23971 23634 23974
rect 23614 23799 23628 23971
rect 23752 23901 23766 24345
rect 24114 24340 24140 24343
rect 24114 24311 24140 24314
rect 23930 24272 23956 24275
rect 23930 24243 23956 24246
rect 23746 23898 23772 23901
rect 23746 23869 23772 23872
rect 23936 23867 23950 24243
rect 24120 24071 24134 24311
rect 24620 24306 24646 24309
rect 24620 24277 24646 24280
rect 24436 24136 24462 24139
rect 24436 24107 24462 24110
rect 24252 24102 24278 24105
rect 24252 24073 24278 24076
rect 24114 24068 24140 24071
rect 24114 24039 24140 24042
rect 24120 24003 24134 24039
rect 24114 24000 24140 24003
rect 24114 23971 24140 23974
rect 23930 23864 23956 23867
rect 23930 23835 23956 23838
rect 23608 23796 23634 23799
rect 23608 23767 23634 23770
rect 23614 23595 23628 23767
rect 23384 23555 23444 23569
rect 23608 23592 23634 23595
rect 23608 23563 23634 23566
rect 23384 23459 23398 23555
rect 23424 23524 23450 23527
rect 23424 23495 23450 23498
rect 24120 23501 24134 23971
rect 24258 23901 24272 24073
rect 24252 23898 24278 23901
rect 24252 23869 24278 23872
rect 23378 23456 23404 23459
rect 23378 23427 23404 23430
rect 23378 22912 23404 22915
rect 23378 22883 23404 22886
rect 23286 22742 23312 22745
rect 23286 22713 23312 22716
rect 23292 22541 23306 22713
rect 23332 22640 23358 22643
rect 23332 22611 23358 22614
rect 23286 22538 23312 22541
rect 23286 22509 23312 22512
rect 23338 22507 23352 22611
rect 23332 22504 23358 22507
rect 23332 22475 23358 22478
rect 23338 22201 23352 22475
rect 23384 22439 23398 22883
rect 23378 22436 23404 22439
rect 23378 22407 23404 22410
rect 23332 22198 23358 22201
rect 23358 22178 23398 22192
rect 23332 22169 23358 22172
rect 23240 21892 23266 21895
rect 23240 21863 23266 21866
rect 23332 21892 23358 21895
rect 23332 21863 23358 21866
rect 23194 21858 23220 21861
rect 23194 21829 23220 21832
rect 23056 20532 23082 20535
rect 23056 20503 23082 20506
rect 23062 20025 23076 20503
rect 23240 20464 23266 20467
rect 23240 20435 23266 20438
rect 23056 20022 23082 20025
rect 23056 19993 23082 19996
rect 23148 20022 23174 20025
rect 23174 20002 23214 20016
rect 23148 19993 23174 19996
rect 23062 19447 23076 19993
rect 23102 19920 23128 19923
rect 23102 19891 23128 19894
rect 23056 19444 23082 19447
rect 23056 19415 23082 19418
rect 23108 19379 23122 19891
rect 23200 19481 23214 20002
rect 23194 19478 23220 19481
rect 23194 19449 23220 19452
rect 23102 19376 23128 19379
rect 23102 19347 23128 19350
rect 23200 18937 23214 19449
rect 23246 18937 23260 20435
rect 23286 20192 23312 20195
rect 23286 20163 23312 20166
rect 23292 20059 23306 20163
rect 23286 20056 23312 20059
rect 23286 20027 23312 20030
rect 23292 19719 23306 20027
rect 23286 19716 23312 19719
rect 23286 19687 23312 19690
rect 23194 18934 23220 18937
rect 23154 18914 23194 18928
rect 23154 18597 23168 18914
rect 23194 18905 23220 18908
rect 23240 18934 23266 18937
rect 23240 18905 23266 18908
rect 23148 18594 23174 18597
rect 23148 18565 23174 18568
rect 23055 18476 23083 18480
rect 23055 18443 23083 18448
rect 23062 18427 23076 18443
rect 23056 18424 23082 18427
rect 23056 18395 23082 18398
rect 23062 18189 23076 18395
rect 23154 18393 23168 18565
rect 23148 18390 23174 18393
rect 23148 18361 23174 18364
rect 23148 18288 23174 18291
rect 23148 18259 23174 18262
rect 23056 18186 23082 18189
rect 23056 18157 23082 18160
rect 23154 17747 23168 18259
rect 23246 18121 23260 18905
rect 23240 18118 23266 18121
rect 23240 18089 23266 18092
rect 23148 17744 23174 17747
rect 23148 17715 23174 17718
rect 23102 17540 23128 17543
rect 23102 17511 23128 17514
rect 23108 17305 23122 17511
rect 23102 17302 23128 17305
rect 23102 17273 23128 17276
rect 23010 16826 23036 16829
rect 23010 16797 23036 16800
rect 23108 16761 23122 17273
rect 23154 17203 23168 17715
rect 23239 17388 23267 17392
rect 23239 17355 23267 17360
rect 23246 17339 23260 17355
rect 23240 17336 23266 17339
rect 23240 17307 23266 17310
rect 23148 17200 23174 17203
rect 23148 17171 23174 17174
rect 23102 16758 23128 16761
rect 23102 16729 23128 16732
rect 23154 16659 23168 17171
rect 23148 16656 23174 16659
rect 23148 16627 23174 16630
rect 23154 16115 23168 16627
rect 23148 16112 23174 16115
rect 23148 16083 23174 16086
rect 22964 15840 22990 15843
rect 22964 15811 22990 15814
rect 22872 15364 22898 15367
rect 22872 15335 22898 15338
rect 22918 15364 22944 15367
rect 22918 15335 22944 15338
rect 22872 15296 22898 15299
rect 22872 15267 22898 15270
rect 22878 14279 22892 15267
rect 22924 14483 22938 15335
rect 22970 15333 22984 15811
rect 22964 15330 22990 15333
rect 22964 15301 22990 15304
rect 22918 14480 22944 14483
rect 22918 14451 22944 14454
rect 22872 14276 22898 14279
rect 22872 14247 22898 14250
rect 22826 14106 22852 14109
rect 22826 14077 22852 14080
rect 22832 13191 22846 14077
rect 22924 13939 22938 14451
rect 23102 14242 23128 14245
rect 23102 14213 23128 14216
rect 22918 13936 22944 13939
rect 22918 13907 22944 13910
rect 23108 13735 23122 14213
rect 23102 13732 23128 13735
rect 23102 13703 23128 13706
rect 23148 13732 23174 13735
rect 23148 13703 23174 13706
rect 23154 13259 23168 13703
rect 23148 13256 23174 13259
rect 23148 13227 23174 13230
rect 22826 13188 22852 13191
rect 22826 13159 22852 13162
rect 22780 13018 22806 13021
rect 22780 12989 22806 12992
rect 22832 12987 22846 13159
rect 22872 13120 22898 13123
rect 22872 13091 22898 13094
rect 22826 12984 22852 12987
rect 22826 12955 22852 12958
rect 22878 12885 22892 13091
rect 22918 12950 22944 12953
rect 22918 12921 22944 12924
rect 22872 12882 22898 12885
rect 22872 12853 22898 12856
rect 22924 11049 22938 12921
rect 22694 11033 22754 11047
rect 22918 11046 22944 11049
rect 23338 11047 23352 21863
rect 23384 21079 23398 22178
rect 23378 21076 23404 21079
rect 23378 21047 23404 21050
rect 23384 20535 23398 21047
rect 23378 20532 23404 20535
rect 23378 20503 23404 20506
rect 23430 18265 23444 23495
rect 24120 23487 24180 23501
rect 24166 22711 24180 23487
rect 24258 22711 24272 23869
rect 24390 23830 24416 23833
rect 24390 23801 24416 23804
rect 24396 23493 24410 23801
rect 24442 23527 24456 24107
rect 24626 24071 24640 24277
rect 24620 24068 24646 24071
rect 24620 24039 24646 24042
rect 24804 24034 24830 24037
rect 24804 24005 24830 24008
rect 24528 23728 24554 23731
rect 24528 23699 24554 23702
rect 24436 23524 24462 23527
rect 24436 23495 24462 23498
rect 24390 23490 24416 23493
rect 24390 23461 24416 23464
rect 24396 22983 24410 23461
rect 24390 22980 24416 22983
rect 24390 22951 24416 22954
rect 24160 22708 24186 22711
rect 24252 22708 24278 22711
rect 24186 22682 24226 22685
rect 24160 22679 24226 22682
rect 24278 22682 24318 22685
rect 24252 22679 24318 22682
rect 24166 22671 24226 22679
rect 24258 22671 24318 22679
rect 24212 22167 24226 22671
rect 24252 22640 24278 22643
rect 24252 22611 24278 22614
rect 24258 22473 24272 22611
rect 24252 22470 24278 22473
rect 24252 22441 24278 22444
rect 24304 22167 24318 22671
rect 24396 22473 24410 22951
rect 24534 22949 24548 23699
rect 24810 23459 24824 24005
rect 24804 23456 24830 23459
rect 24804 23427 24830 23430
rect 24528 22946 24554 22949
rect 24528 22917 24554 22920
rect 24390 22470 24416 22473
rect 24390 22441 24416 22444
rect 24344 22402 24370 22405
rect 24344 22373 24370 22376
rect 24350 22235 24364 22373
rect 24344 22232 24370 22235
rect 24344 22203 24370 22206
rect 24206 22164 24232 22167
rect 24206 22135 24232 22138
rect 24298 22164 24324 22167
rect 24298 22135 24324 22138
rect 23700 21382 23726 21385
rect 23700 21353 23726 21356
rect 23706 21113 23720 21353
rect 23884 21178 23910 21181
rect 23884 21149 23910 21152
rect 23700 21110 23726 21113
rect 23700 21081 23726 21084
rect 23562 20566 23588 20569
rect 23562 20537 23588 20540
rect 23654 20566 23680 20569
rect 23706 20560 23720 21081
rect 23890 21011 23904 21149
rect 23884 21008 23910 21011
rect 23884 20979 23910 20982
rect 23890 20707 23904 20979
rect 23890 20693 23950 20707
rect 23936 20569 23950 20693
rect 23680 20546 23720 20560
rect 23930 20566 23956 20569
rect 23654 20537 23680 20540
rect 23930 20537 23956 20540
rect 23568 20025 23582 20537
rect 24114 20192 24140 20195
rect 24114 20163 24140 20166
rect 24120 20059 24134 20163
rect 24114 20056 24140 20059
rect 24114 20027 24140 20030
rect 23562 20022 23588 20025
rect 23562 19993 23588 19996
rect 24160 19104 24186 19107
rect 24160 19075 24186 19078
rect 24114 18968 24140 18971
rect 24114 18939 24140 18942
rect 24022 18866 24048 18869
rect 24022 18837 24048 18840
rect 22694 11015 22708 11033
rect 22878 11026 22918 11040
rect 22688 11012 22714 11015
rect 22688 10983 22714 10986
rect 22596 10978 22622 10981
rect 22596 10949 22622 10952
rect 22642 10978 22668 10981
rect 22642 10949 22668 10952
rect 22550 9890 22576 9893
rect 22550 9861 22576 9864
rect 22556 9689 22570 9861
rect 22550 9686 22576 9689
rect 22550 9657 22576 9660
rect 22556 9417 22570 9657
rect 22550 9414 22576 9417
rect 22550 9385 22576 9388
rect 22411 9364 22439 9368
rect 22411 9331 22439 9336
rect 22602 9213 22616 10949
rect 22648 10845 22662 10949
rect 22642 10842 22668 10845
rect 22642 10813 22668 10816
rect 22694 10456 22708 10983
rect 22687 10452 22715 10456
rect 22687 10419 22715 10424
rect 22826 10298 22852 10301
rect 22826 10269 22852 10272
rect 22642 9958 22668 9961
rect 22642 9929 22668 9932
rect 22648 9723 22662 9929
rect 22688 9924 22714 9927
rect 22688 9895 22714 9898
rect 22642 9720 22668 9723
rect 22642 9691 22668 9694
rect 22648 9383 22662 9691
rect 22694 9689 22708 9895
rect 22734 9890 22760 9893
rect 22734 9861 22760 9864
rect 22740 9689 22754 9861
rect 22688 9686 22714 9689
rect 22688 9657 22714 9660
rect 22734 9686 22760 9689
rect 22734 9657 22760 9660
rect 22694 9383 22708 9657
rect 22642 9380 22668 9383
rect 22642 9351 22668 9354
rect 22688 9380 22714 9383
rect 22688 9351 22714 9354
rect 22596 9210 22622 9213
rect 22596 9181 22622 9184
rect 22648 9145 22662 9351
rect 22642 9142 22668 9145
rect 22642 9113 22668 9116
rect 22648 8873 22662 9113
rect 22694 9077 22708 9351
rect 22740 9179 22754 9657
rect 22780 9414 22806 9417
rect 22780 9385 22806 9388
rect 22734 9176 22760 9179
rect 22734 9147 22760 9150
rect 22786 9145 22800 9385
rect 22780 9142 22806 9145
rect 22780 9113 22806 9116
rect 22688 9074 22714 9077
rect 22688 9045 22714 9048
rect 22642 8870 22668 8873
rect 22642 8841 22668 8844
rect 22596 8802 22622 8805
rect 22596 8773 22622 8776
rect 22602 8601 22616 8773
rect 22648 8601 22662 8841
rect 22694 8805 22708 9045
rect 22786 8839 22800 9113
rect 22780 8836 22806 8839
rect 22780 8807 22806 8810
rect 22688 8802 22714 8805
rect 22688 8773 22714 8776
rect 22734 8768 22760 8771
rect 22734 8739 22760 8742
rect 22596 8598 22622 8601
rect 22596 8569 22622 8572
rect 22642 8598 22668 8601
rect 22642 8569 22668 8572
rect 22648 8329 22662 8569
rect 22688 8530 22714 8533
rect 22688 8501 22714 8504
rect 22642 8326 22668 8329
rect 22642 8297 22668 8300
rect 22694 8295 22708 8501
rect 22688 8292 22714 8295
rect 22688 8263 22714 8266
rect 22694 7751 22708 8263
rect 22740 8125 22754 8739
rect 22786 8601 22800 8807
rect 22780 8598 22806 8601
rect 22780 8569 22806 8572
rect 22786 8295 22800 8569
rect 22780 8292 22806 8295
rect 22780 8263 22806 8266
rect 22734 8122 22760 8125
rect 22734 8093 22760 8096
rect 22688 7748 22714 7751
rect 22648 7728 22688 7742
rect 22648 7207 22662 7728
rect 22688 7719 22714 7722
rect 22688 7476 22714 7479
rect 22688 7447 22714 7450
rect 22642 7204 22668 7207
rect 22642 7175 22668 7178
rect 22596 7136 22622 7139
rect 22596 7107 22622 7110
rect 22602 6969 22616 7107
rect 22596 6966 22622 6969
rect 22596 6937 22622 6940
rect 22642 6966 22668 6969
rect 22642 6937 22668 6940
rect 22602 6920 22616 6937
rect 22595 6916 22623 6920
rect 22595 6883 22623 6888
rect 22648 6765 22662 6937
rect 22642 6762 22668 6765
rect 22642 6733 22668 6736
rect 22694 5575 22708 7447
rect 22740 7028 22754 8093
rect 22786 7785 22800 8263
rect 22832 8227 22846 10269
rect 22878 8669 22892 11026
rect 22918 11017 22944 11020
rect 23108 11033 23352 11047
rect 23384 18251 23444 18265
rect 23010 10978 23036 10981
rect 23010 10949 23036 10952
rect 22917 10792 22945 10796
rect 22917 10759 22918 10764
rect 22944 10759 22945 10764
rect 22918 10745 22944 10748
rect 23016 10573 23030 10949
rect 23108 10777 23122 11033
rect 23148 11012 23174 11015
rect 23148 10983 23174 10986
rect 23240 11012 23266 11015
rect 23240 10983 23266 10986
rect 23102 10774 23128 10777
rect 23102 10745 23128 10748
rect 23010 10570 23036 10573
rect 23010 10541 23036 10544
rect 23108 10471 23122 10745
rect 23154 10573 23168 10983
rect 23194 10944 23220 10947
rect 23194 10915 23220 10918
rect 23200 10811 23214 10915
rect 23246 10845 23260 10983
rect 23240 10842 23266 10845
rect 23240 10813 23266 10816
rect 23194 10808 23220 10811
rect 23384 10796 23398 18251
rect 23424 18118 23450 18121
rect 23424 18089 23450 18092
rect 23194 10779 23220 10782
rect 23377 10792 23405 10796
rect 23377 10759 23405 10764
rect 23240 10740 23266 10743
rect 23430 10717 23444 18089
rect 23976 17846 24002 17849
rect 23976 17817 24002 17820
rect 23982 17611 23996 17817
rect 23976 17608 24002 17611
rect 23976 17579 24002 17582
rect 23982 17528 23996 17579
rect 23975 17524 24003 17528
rect 23975 17491 24003 17496
rect 24028 16557 24042 18837
rect 24120 18665 24134 18939
rect 24114 18662 24140 18665
rect 24114 18633 24140 18636
rect 24166 18631 24180 19075
rect 24160 18628 24186 18631
rect 24160 18599 24186 18602
rect 24166 18291 24180 18599
rect 24160 18288 24186 18291
rect 24160 18259 24186 18262
rect 24068 17846 24094 17849
rect 24068 17817 24094 17820
rect 24074 17645 24088 17817
rect 24068 17642 24094 17645
rect 24068 17613 24094 17616
rect 24166 17543 24180 18259
rect 24160 17540 24186 17543
rect 24160 17511 24186 17514
rect 24114 16656 24140 16659
rect 24114 16627 24140 16630
rect 24022 16554 24048 16557
rect 24022 16525 24048 16528
rect 24120 16455 24134 16627
rect 24114 16452 24140 16455
rect 24114 16423 24140 16426
rect 23976 16418 24002 16421
rect 23976 16389 24002 16392
rect 23982 16285 23996 16389
rect 23976 16282 24002 16285
rect 23976 16253 24002 16256
rect 24160 15908 24186 15911
rect 24160 15879 24186 15882
rect 24166 15401 24180 15879
rect 24160 15398 24186 15401
rect 24160 15369 24186 15372
rect 24166 14857 24180 15369
rect 24160 14854 24186 14857
rect 24160 14825 24186 14828
rect 24114 14106 24140 14109
rect 24114 14077 24140 14080
rect 24068 13800 24094 13803
rect 24068 13771 24094 13774
rect 23929 12968 23957 12972
rect 23929 12935 23957 12940
rect 23936 12307 23950 12935
rect 24074 12375 24088 13771
rect 24068 12372 24094 12375
rect 24068 12343 24094 12346
rect 23930 12304 23956 12307
rect 23930 12275 23956 12278
rect 23976 11012 24002 11015
rect 23976 10983 24002 10986
rect 23515 10860 23543 10864
rect 23515 10827 23516 10832
rect 23542 10827 23543 10832
rect 23516 10813 23542 10816
rect 23240 10711 23266 10714
rect 23246 10675 23260 10711
rect 23384 10703 23444 10717
rect 23240 10672 23266 10675
rect 23240 10643 23266 10646
rect 23148 10570 23174 10573
rect 23148 10541 23174 10544
rect 23102 10468 23128 10471
rect 23102 10439 23128 10442
rect 23108 9995 23122 10439
rect 23102 9992 23128 9995
rect 23102 9963 23128 9966
rect 23246 9417 23260 10643
rect 23240 9414 23266 9417
rect 23240 9385 23266 9388
rect 22963 9364 22991 9368
rect 22963 9331 22991 9336
rect 22970 9315 22984 9331
rect 22964 9312 22990 9315
rect 22964 9283 22990 9286
rect 22872 8666 22898 8669
rect 22872 8637 22898 8640
rect 23246 8601 23260 9385
rect 23384 9153 23398 10703
rect 23562 10672 23588 10675
rect 23522 10652 23562 10666
rect 23522 10471 23536 10652
rect 23562 10643 23588 10646
rect 23982 10573 23996 10983
rect 24022 10944 24048 10947
rect 24022 10915 24048 10918
rect 24028 10811 24042 10915
rect 24022 10808 24048 10811
rect 24022 10779 24048 10782
rect 24120 10573 24134 14077
rect 24160 13460 24186 13463
rect 24160 13431 24186 13434
rect 24166 13293 24180 13431
rect 24160 13290 24186 13293
rect 24160 13261 24186 13264
rect 24212 11047 24226 22135
rect 24396 21929 24410 22441
rect 24534 22439 24548 22917
rect 24528 22436 24554 22439
rect 24488 22410 24528 22413
rect 24488 22407 24554 22410
rect 24436 22402 24462 22405
rect 24436 22373 24462 22376
rect 24488 22399 24548 22407
rect 24442 22356 24456 22373
rect 24435 22352 24463 22356
rect 24435 22319 24463 22324
rect 24390 21926 24416 21929
rect 24390 21897 24416 21900
rect 24396 21419 24410 21897
rect 24488 21861 24502 22399
rect 24482 21858 24508 21861
rect 24482 21829 24508 21832
rect 24666 21858 24692 21861
rect 24666 21829 24692 21832
rect 24390 21416 24416 21419
rect 24390 21387 24416 21390
rect 24488 21385 24502 21829
rect 24672 21691 24686 21829
rect 24666 21688 24692 21691
rect 24666 21659 24692 21662
rect 24482 21382 24508 21385
rect 24482 21353 24508 21356
rect 24620 21348 24646 21351
rect 24620 21319 24646 21322
rect 24574 21008 24600 21011
rect 24574 20979 24600 20982
rect 24580 20773 24594 20979
rect 24626 20773 24640 21319
rect 24758 21314 24784 21317
rect 24758 21285 24784 21288
rect 24666 20838 24692 20841
rect 24666 20809 24692 20812
rect 24574 20770 24600 20773
rect 24574 20741 24600 20744
rect 24620 20770 24646 20773
rect 24620 20741 24646 20744
rect 24436 20022 24462 20025
rect 24436 19993 24462 19996
rect 24482 20022 24508 20025
rect 24482 19993 24508 19996
rect 24252 19920 24278 19923
rect 24252 19891 24278 19894
rect 24298 19920 24324 19923
rect 24298 19891 24324 19894
rect 24258 19821 24272 19891
rect 24252 19818 24278 19821
rect 24252 19789 24278 19792
rect 24304 19005 24318 19891
rect 24389 19564 24417 19568
rect 24442 19549 24456 19993
rect 24488 19923 24502 19993
rect 24482 19920 24508 19923
rect 24482 19891 24508 19894
rect 24488 19787 24502 19891
rect 24482 19784 24508 19787
rect 24482 19755 24508 19758
rect 24389 19531 24417 19536
rect 24436 19546 24462 19549
rect 24298 19002 24324 19005
rect 24298 18973 24324 18976
rect 24252 18934 24278 18937
rect 24252 18905 24278 18908
rect 24344 18934 24370 18937
rect 24344 18905 24370 18908
rect 24258 17917 24272 18905
rect 24298 18832 24324 18835
rect 24298 18803 24324 18806
rect 24304 18427 24318 18803
rect 24298 18424 24324 18427
rect 24298 18395 24324 18398
rect 24350 18359 24364 18905
rect 24396 18393 24410 19531
rect 24436 19517 24462 19520
rect 24436 19138 24462 19141
rect 24436 19109 24462 19112
rect 24442 18971 24456 19109
rect 24672 19005 24686 20809
rect 24764 20807 24778 21285
rect 24758 20804 24784 20807
rect 24758 20775 24784 20778
rect 24712 20770 24738 20773
rect 24712 20741 24738 20744
rect 24718 20637 24732 20741
rect 24712 20634 24738 20637
rect 24712 20605 24738 20608
rect 24666 19002 24692 19005
rect 24666 18973 24692 18976
rect 24436 18968 24462 18971
rect 24436 18939 24462 18942
rect 24666 18832 24692 18835
rect 24666 18803 24692 18806
rect 24481 18612 24509 18616
rect 24481 18579 24482 18584
rect 24508 18579 24509 18584
rect 24482 18565 24508 18568
rect 24481 18408 24509 18412
rect 24390 18390 24416 18393
rect 24481 18375 24482 18380
rect 24390 18361 24416 18364
rect 24508 18375 24509 18380
rect 24482 18361 24508 18364
rect 24344 18356 24370 18359
rect 24344 18327 24370 18330
rect 24482 18322 24508 18325
rect 24482 18293 24508 18296
rect 24252 17914 24278 17917
rect 24252 17885 24278 17888
rect 24298 17778 24324 17781
rect 24298 17749 24324 17752
rect 24304 17237 24318 17749
rect 24436 17540 24462 17543
rect 24436 17511 24462 17514
rect 24298 17234 24324 17237
rect 24298 17205 24324 17208
rect 24442 17101 24456 17511
rect 24436 17098 24462 17101
rect 24436 17069 24462 17072
rect 24390 15874 24416 15877
rect 24390 15845 24416 15848
rect 24396 15707 24410 15845
rect 24390 15704 24416 15707
rect 24390 15675 24416 15678
rect 24396 15367 24410 15675
rect 24390 15364 24416 15367
rect 24390 15335 24416 15338
rect 24344 14854 24370 14857
rect 24344 14825 24370 14828
rect 24298 14480 24324 14483
rect 24298 14451 24324 14454
rect 24252 13392 24278 13395
rect 24252 13363 24278 13366
rect 24258 12477 24272 13363
rect 24252 12474 24278 12477
rect 24252 12445 24278 12448
rect 24304 11321 24318 14451
rect 24350 14313 24364 14825
rect 24390 14820 24416 14823
rect 24390 14791 24416 14794
rect 24344 14310 24370 14313
rect 24344 14281 24370 14284
rect 24350 13769 24364 14281
rect 24396 14245 24410 14791
rect 24390 14242 24416 14245
rect 24390 14213 24416 14216
rect 24396 14041 24410 14213
rect 24390 14038 24416 14041
rect 24390 14009 24416 14012
rect 24344 13766 24370 13769
rect 24344 13737 24370 13740
rect 24396 13735 24410 14009
rect 24390 13732 24416 13735
rect 24390 13703 24416 13706
rect 24436 12406 24462 12409
rect 24436 12377 24462 12380
rect 24442 11389 24456 12377
rect 24436 11386 24462 11389
rect 24436 11357 24462 11360
rect 24298 11318 24324 11321
rect 24298 11289 24324 11292
rect 24166 11033 24226 11047
rect 23976 10570 24002 10573
rect 23976 10541 24002 10544
rect 24114 10570 24140 10573
rect 24114 10541 24140 10544
rect 23516 10468 23542 10471
rect 23423 10452 23451 10456
rect 23516 10439 23542 10442
rect 23423 10419 23451 10424
rect 23430 9757 23444 10419
rect 23424 9754 23450 9757
rect 23424 9725 23450 9728
rect 23424 9380 23450 9383
rect 23424 9351 23450 9354
rect 23430 9213 23444 9351
rect 23424 9210 23450 9213
rect 23424 9181 23450 9184
rect 23384 9139 23444 9153
rect 23522 9145 23536 10439
rect 24120 10301 24134 10541
rect 24166 10403 24180 11033
rect 24160 10400 24186 10403
rect 24160 10371 24186 10374
rect 24114 10298 24140 10301
rect 24114 10269 24140 10272
rect 23976 9482 24002 9485
rect 23976 9453 24002 9456
rect 23884 9448 23910 9451
rect 23884 9419 23910 9422
rect 23838 9414 23864 9417
rect 23838 9385 23864 9388
rect 23240 8598 23266 8601
rect 23240 8569 23266 8572
rect 22964 8564 22990 8567
rect 22964 8535 22990 8538
rect 22970 8295 22984 8535
rect 22964 8292 22990 8295
rect 22964 8263 22990 8266
rect 22918 8258 22944 8261
rect 22918 8229 22944 8232
rect 22826 8224 22852 8227
rect 22826 8195 22852 8198
rect 22780 7782 22806 7785
rect 22780 7753 22806 7756
rect 22786 7207 22800 7753
rect 22780 7204 22806 7207
rect 22780 7175 22806 7178
rect 22924 7139 22938 8229
rect 22964 8224 22990 8227
rect 22964 8195 22990 8198
rect 23010 8224 23036 8227
rect 23010 8195 23036 8198
rect 22918 7136 22944 7139
rect 22918 7107 22944 7110
rect 22740 7014 22800 7028
rect 22734 6966 22760 6969
rect 22734 6937 22760 6940
rect 22740 6493 22754 6937
rect 22786 6901 22800 7014
rect 22924 6969 22938 7107
rect 22918 6966 22944 6969
rect 22918 6937 22944 6940
rect 22780 6898 22806 6901
rect 22780 6869 22806 6872
rect 22734 6490 22760 6493
rect 22734 6461 22760 6464
rect 22970 6323 22984 8195
rect 23016 8125 23030 8195
rect 23010 8122 23036 8125
rect 23010 8093 23036 8096
rect 23246 8057 23260 8569
rect 23430 8091 23444 9139
rect 23516 9142 23542 9145
rect 23516 9113 23542 9116
rect 23522 8601 23536 9113
rect 23844 9111 23858 9385
rect 23890 9179 23904 9419
rect 23982 9315 23996 9453
rect 24206 9346 24232 9349
rect 24206 9317 24232 9320
rect 23976 9312 24002 9315
rect 23976 9283 24002 9286
rect 23884 9176 23910 9179
rect 23883 9160 23884 9164
rect 23910 9160 23911 9164
rect 23982 9145 23996 9283
rect 23883 9127 23911 9132
rect 23976 9142 24002 9145
rect 23976 9113 24002 9116
rect 23838 9108 23864 9111
rect 23838 9079 23864 9082
rect 24212 9043 24226 9317
rect 24206 9040 24232 9043
rect 24205 9024 24206 9028
rect 24232 9024 24233 9028
rect 24205 8991 24233 8996
rect 23608 8768 23634 8771
rect 23608 8739 23634 8742
rect 23614 8635 23628 8739
rect 23608 8632 23634 8635
rect 23608 8603 23634 8606
rect 23516 8598 23542 8601
rect 23516 8569 23542 8572
rect 23424 8088 23450 8091
rect 23424 8059 23450 8062
rect 23240 8054 23266 8057
rect 23240 8025 23266 8028
rect 23246 7513 23260 8025
rect 23240 7510 23266 7513
rect 23240 7481 23266 7484
rect 23246 7309 23260 7481
rect 23240 7306 23266 7309
rect 23240 7277 23266 7280
rect 23246 6969 23260 7277
rect 23240 6966 23266 6969
rect 23240 6937 23266 6940
rect 23246 6697 23260 6937
rect 23240 6694 23266 6697
rect 23240 6665 23266 6668
rect 23246 6433 23260 6665
rect 23430 6512 23444 8059
rect 23522 8057 23536 8569
rect 24344 8496 24370 8499
rect 24344 8467 24370 8470
rect 24298 8360 24324 8363
rect 24298 8331 24324 8334
rect 24304 8227 24318 8331
rect 24350 8295 24364 8467
rect 24488 8397 24502 18293
rect 24620 17540 24646 17543
rect 24620 17511 24646 17514
rect 24528 17506 24554 17509
rect 24528 17477 24554 17480
rect 24534 16217 24548 17477
rect 24574 16996 24600 16999
rect 24626 16990 24640 17511
rect 24600 16976 24640 16990
rect 24574 16967 24600 16970
rect 24528 16214 24554 16217
rect 24528 16185 24554 16188
rect 24534 15877 24548 16185
rect 24534 15874 24600 15877
rect 24534 15863 24574 15874
rect 24574 15845 24600 15848
rect 24580 14245 24594 15845
rect 24672 14279 24686 18803
rect 24712 17268 24738 17271
rect 24712 17239 24738 17242
rect 24718 17101 24732 17239
rect 24712 17098 24738 17101
rect 24712 17069 24738 17072
rect 24712 16520 24738 16523
rect 24712 16491 24738 16494
rect 24666 14276 24692 14279
rect 24666 14247 24692 14250
rect 24574 14242 24600 14245
rect 24574 14213 24600 14216
rect 24718 13701 24732 16491
rect 24810 15877 24824 23427
rect 24850 22946 24876 22949
rect 24850 22917 24876 22920
rect 24856 22779 24870 22917
rect 25632 22912 25658 22915
rect 25632 22883 25658 22886
rect 24850 22776 24876 22779
rect 24850 22747 24876 22750
rect 25402 22368 25428 22371
rect 25402 22339 25428 22342
rect 25408 22201 25422 22339
rect 25638 22235 25652 22883
rect 28254 22776 28280 22779
rect 28254 22747 28280 22750
rect 28208 22708 28234 22711
rect 28208 22679 28234 22682
rect 26966 22436 26992 22439
rect 26966 22407 26992 22410
rect 25632 22232 25658 22235
rect 25632 22203 25658 22206
rect 26230 22232 26256 22235
rect 26230 22203 26256 22206
rect 25402 22198 25428 22201
rect 25402 22169 25428 22172
rect 25586 22198 25612 22201
rect 25586 22169 25612 22172
rect 25592 21997 25606 22169
rect 26138 22164 26164 22167
rect 26138 22135 26164 22138
rect 25678 22096 25704 22099
rect 25678 22067 25704 22070
rect 25586 21994 25612 21997
rect 25586 21965 25612 21968
rect 25632 21960 25658 21963
rect 25632 21931 25658 21934
rect 25540 21620 25566 21623
rect 25540 21591 25566 21594
rect 25546 21419 25560 21591
rect 25540 21416 25566 21419
rect 25540 21387 25566 21390
rect 25546 21113 25560 21387
rect 25540 21110 25566 21113
rect 25540 21081 25566 21084
rect 25546 20535 25560 21081
rect 25586 20600 25612 20603
rect 25586 20571 25612 20574
rect 25540 20532 25566 20535
rect 25540 20503 25566 20506
rect 25546 20025 25560 20503
rect 25592 20365 25606 20571
rect 25586 20362 25612 20365
rect 25586 20333 25612 20336
rect 25540 20022 25566 20025
rect 25540 19993 25566 19996
rect 25540 19274 25566 19277
rect 25540 19245 25566 19248
rect 25494 19104 25520 19107
rect 25494 19075 25520 19078
rect 25500 18971 25514 19075
rect 25494 18968 25520 18971
rect 25494 18939 25520 18942
rect 25356 18934 25382 18937
rect 25356 18905 25382 18908
rect 25448 18934 25474 18937
rect 25448 18905 25474 18908
rect 25362 18733 25376 18905
rect 25356 18730 25382 18733
rect 25356 18701 25382 18704
rect 25454 18699 25468 18905
rect 25546 18877 25560 19245
rect 25500 18869 25560 18877
rect 25494 18866 25560 18869
rect 25520 18863 25560 18866
rect 25494 18837 25520 18840
rect 25448 18696 25474 18699
rect 25448 18667 25474 18670
rect 25592 17392 25606 20333
rect 25638 19277 25652 21931
rect 25684 21895 25698 22067
rect 26144 21895 26158 22135
rect 26184 21994 26210 21997
rect 26184 21965 26210 21968
rect 25678 21892 25704 21895
rect 25862 21892 25888 21895
rect 25678 21863 25704 21866
rect 25861 21876 25862 21880
rect 26138 21892 26164 21895
rect 25888 21876 25889 21880
rect 26138 21863 26164 21866
rect 25861 21843 25889 21848
rect 25868 21725 25882 21843
rect 25862 21722 25888 21725
rect 25862 21693 25888 21696
rect 26144 21623 26158 21863
rect 26138 21620 26164 21623
rect 26138 21591 26164 21594
rect 26190 21453 26204 21965
rect 26236 21929 26250 22203
rect 26874 22198 26900 22201
rect 26874 22169 26900 22172
rect 26230 21926 26256 21929
rect 26230 21897 26256 21900
rect 26880 21895 26894 22169
rect 26874 21892 26900 21895
rect 26874 21863 26900 21866
rect 26368 21688 26394 21691
rect 26368 21659 26394 21662
rect 26184 21450 26210 21453
rect 26184 21421 26210 21424
rect 25724 21076 25750 21079
rect 25724 21047 25750 21050
rect 25730 20707 25744 21047
rect 26374 21011 26388 21659
rect 26880 21657 26894 21863
rect 26972 21861 26986 22407
rect 28214 22201 28228 22679
rect 28208 22198 28234 22201
rect 28208 22169 28234 22172
rect 27150 22096 27176 22099
rect 27150 22067 27176 22070
rect 28024 22096 28050 22099
rect 28024 22067 28050 22070
rect 27156 21948 27170 22067
rect 27380 21994 27406 21997
rect 27380 21965 27406 21968
rect 27149 21944 27177 21948
rect 27110 21923 27149 21937
rect 26966 21858 26992 21861
rect 26966 21829 26992 21832
rect 26874 21654 26900 21657
rect 26874 21625 26900 21628
rect 26880 21113 26894 21625
rect 26874 21110 26900 21113
rect 26874 21081 26900 21084
rect 26368 21008 26394 21011
rect 26368 20979 26394 20982
rect 26880 20841 26894 21081
rect 27012 21008 27038 21011
rect 27012 20979 27038 20982
rect 26874 20838 26900 20841
rect 26874 20809 26900 20812
rect 25684 20693 25744 20707
rect 25684 20569 25698 20693
rect 25678 20566 25704 20569
rect 25678 20537 25704 20540
rect 25730 20025 25744 20693
rect 26828 20566 26854 20569
rect 26828 20537 26854 20540
rect 26230 20464 26256 20467
rect 26230 20435 26256 20438
rect 26782 20464 26808 20467
rect 26782 20435 26808 20438
rect 25724 20022 25750 20025
rect 25724 19993 25750 19996
rect 25632 19274 25658 19277
rect 25632 19245 25658 19248
rect 25730 18937 25744 19993
rect 25632 18934 25658 18937
rect 25632 18905 25658 18908
rect 25724 18934 25750 18937
rect 25724 18905 25750 18908
rect 25638 17543 25652 18905
rect 26236 18665 26250 20435
rect 26788 20263 26802 20435
rect 26834 20365 26848 20537
rect 26828 20362 26854 20365
rect 26828 20333 26854 20336
rect 27018 20331 27032 20979
rect 27058 20804 27084 20807
rect 27058 20775 27084 20778
rect 27012 20328 27038 20331
rect 27012 20299 27038 20302
rect 27064 20263 27078 20775
rect 26322 20260 26348 20263
rect 26322 20231 26348 20234
rect 26782 20260 26808 20263
rect 26782 20231 26808 20234
rect 27058 20260 27084 20263
rect 27058 20231 27084 20234
rect 26230 18662 26256 18665
rect 26230 18633 26256 18636
rect 26230 18594 26256 18597
rect 26230 18565 26256 18568
rect 26276 18594 26302 18597
rect 26276 18565 26302 18568
rect 26138 17846 26164 17849
rect 26138 17817 26164 17820
rect 25724 17744 25750 17747
rect 25724 17715 25750 17718
rect 25632 17540 25658 17543
rect 25632 17511 25658 17514
rect 25585 17388 25613 17392
rect 25585 17355 25613 17360
rect 25586 17336 25612 17339
rect 25586 17307 25612 17310
rect 25592 16523 25606 17307
rect 25638 17305 25652 17511
rect 25632 17302 25658 17305
rect 25632 17273 25658 17276
rect 25586 16520 25612 16523
rect 25546 16494 25586 16497
rect 25546 16491 25612 16494
rect 25546 16483 25606 16491
rect 25356 16180 25382 16183
rect 25356 16151 25382 16154
rect 25362 15945 25376 16151
rect 25356 15942 25382 15945
rect 25356 15913 25382 15916
rect 24764 15863 24824 15877
rect 24764 14823 24778 15863
rect 25362 15673 25376 15913
rect 25546 15681 25560 16483
rect 25586 15942 25612 15945
rect 25586 15913 25612 15916
rect 25592 15749 25606 15913
rect 25730 15911 25744 17715
rect 26144 17611 26158 17817
rect 26184 17812 26210 17815
rect 26184 17783 26210 17786
rect 26138 17608 26164 17611
rect 26138 17579 26164 17582
rect 26190 17543 26204 17783
rect 25770 17540 25796 17543
rect 25770 17511 25796 17514
rect 26092 17540 26118 17543
rect 26092 17511 26118 17514
rect 26184 17540 26210 17543
rect 26184 17511 26210 17514
rect 25776 17101 25790 17511
rect 25862 17472 25888 17475
rect 25862 17443 25888 17446
rect 25770 17098 25796 17101
rect 25770 17069 25796 17072
rect 25868 16421 25882 17443
rect 25907 17388 25935 17392
rect 25907 17355 25935 17360
rect 25862 16418 25888 16421
rect 25862 16389 25888 16392
rect 25816 15976 25842 15979
rect 25816 15947 25842 15950
rect 25632 15908 25658 15911
rect 25632 15879 25658 15882
rect 25724 15908 25750 15911
rect 25724 15879 25750 15882
rect 25638 15817 25652 15879
rect 25638 15803 25698 15817
rect 25592 15735 25652 15749
rect 25586 15704 25612 15707
rect 25546 15678 25586 15681
rect 25546 15675 25612 15678
rect 25356 15670 25382 15673
rect 25546 15667 25606 15675
rect 25356 15641 25382 15644
rect 24758 14820 24784 14823
rect 24758 14791 24784 14794
rect 25638 14279 25652 15735
rect 25684 15469 25698 15803
rect 25678 15466 25704 15469
rect 25678 15437 25704 15440
rect 25730 15435 25744 15879
rect 25724 15432 25750 15435
rect 25724 15403 25750 15406
rect 25822 14347 25836 15947
rect 25868 15945 25882 16389
rect 25914 16251 25928 17355
rect 26000 16792 26026 16795
rect 26000 16763 26026 16766
rect 25908 16248 25934 16251
rect 25908 16219 25934 16222
rect 25862 15942 25888 15945
rect 25862 15913 25888 15916
rect 25914 15877 25928 16219
rect 25868 15863 25928 15877
rect 25816 14344 25842 14347
rect 25816 14315 25842 14318
rect 25632 14276 25658 14279
rect 25632 14247 25658 14250
rect 25770 14276 25796 14279
rect 25770 14247 25796 14250
rect 25776 13837 25790 14247
rect 25822 14109 25836 14315
rect 25816 14106 25842 14109
rect 25816 14077 25842 14080
rect 25770 13834 25796 13837
rect 25770 13805 25796 13808
rect 25356 13800 25382 13803
rect 25356 13771 25382 13774
rect 24712 13698 24738 13701
rect 24712 13669 24738 13672
rect 24718 13301 24732 13669
rect 25362 13497 25376 13771
rect 25356 13494 25382 13497
rect 25356 13465 25382 13468
rect 24718 13287 24824 13301
rect 24810 12700 24824 13287
rect 25868 12987 25882 15863
rect 26006 15571 26020 16763
rect 26046 16758 26072 16761
rect 26046 16729 26072 16732
rect 26052 16217 26066 16729
rect 26098 16455 26112 17511
rect 26138 17098 26164 17101
rect 26138 17069 26164 17072
rect 26144 16644 26158 17069
rect 26137 16640 26165 16644
rect 26137 16607 26165 16612
rect 26092 16452 26118 16455
rect 26092 16423 26118 16426
rect 26046 16214 26072 16217
rect 26046 16185 26072 16188
rect 26052 15877 26066 16185
rect 26098 15945 26112 16423
rect 26092 15942 26118 15945
rect 26092 15913 26118 15916
rect 26144 15877 26158 16607
rect 26046 15874 26072 15877
rect 26144 15863 26204 15877
rect 26046 15845 26072 15848
rect 26052 15673 26066 15845
rect 26046 15670 26072 15673
rect 26046 15641 26072 15644
rect 26000 15568 26026 15571
rect 26000 15539 26026 15542
rect 25908 14752 25934 14755
rect 25908 14723 25934 14726
rect 25914 14347 25928 14723
rect 26138 14582 26164 14585
rect 26138 14553 26164 14556
rect 26000 14548 26026 14551
rect 26000 14519 26026 14522
rect 25908 14344 25934 14347
rect 25908 14315 25934 14318
rect 26006 14279 26020 14519
rect 26000 14276 26026 14279
rect 26000 14247 26026 14250
rect 25954 14004 25980 14007
rect 26006 13981 26020 14247
rect 26144 14049 26158 14553
rect 26190 14075 26204 15863
rect 26098 14041 26158 14049
rect 26184 14072 26210 14075
rect 26184 14043 26210 14046
rect 26092 14038 26158 14041
rect 26118 14035 26158 14038
rect 26092 14009 26118 14012
rect 25980 13978 26020 13981
rect 25954 13975 26020 13978
rect 25960 13967 26020 13975
rect 26006 13497 26020 13967
rect 26144 13497 26158 14035
rect 26236 13939 26250 18565
rect 26230 13936 26256 13939
rect 26230 13907 26256 13910
rect 26282 13641 26296 18565
rect 26328 17611 26342 20231
rect 26920 20192 26946 20195
rect 26920 20163 26946 20166
rect 26926 20025 26940 20163
rect 26920 20022 26946 20025
rect 26920 19993 26946 19996
rect 26690 19240 26716 19243
rect 26690 19211 26716 19214
rect 26506 18968 26532 18971
rect 26466 18948 26506 18962
rect 26466 18563 26480 18948
rect 26506 18939 26532 18942
rect 26696 18631 26710 19211
rect 27058 18696 27084 18699
rect 27058 18667 27084 18670
rect 26690 18628 26716 18631
rect 26690 18599 26716 18602
rect 26460 18560 26486 18563
rect 26460 18531 26486 18534
rect 26466 17883 26480 18531
rect 26460 17880 26486 17883
rect 26460 17851 26486 17854
rect 26368 17846 26394 17849
rect 26368 17817 26394 17820
rect 26374 17789 26388 17817
rect 26374 17775 26434 17789
rect 26322 17608 26348 17611
rect 26322 17579 26348 17582
rect 26368 17506 26394 17509
rect 26368 17477 26394 17480
rect 26374 17373 26388 17477
rect 26368 17370 26394 17373
rect 26368 17341 26394 17344
rect 26420 16965 26434 17775
rect 26414 16962 26440 16965
rect 26414 16933 26440 16936
rect 26420 16761 26434 16933
rect 26414 16758 26440 16761
rect 26414 16729 26440 16732
rect 26368 15908 26394 15911
rect 26368 15879 26394 15882
rect 26374 15741 26388 15879
rect 26368 15738 26394 15741
rect 26368 15709 26394 15712
rect 26322 15568 26348 15571
rect 26322 15539 26348 15542
rect 26236 13627 26296 13641
rect 26000 13494 26026 13497
rect 26000 13465 26026 13468
rect 26138 13494 26164 13497
rect 26138 13465 26164 13468
rect 25862 12984 25888 12987
rect 25862 12955 25888 12958
rect 25632 12950 25658 12953
rect 25632 12921 25658 12924
rect 25540 12848 25566 12851
rect 25540 12819 25566 12822
rect 24803 12696 24831 12700
rect 24803 12663 24831 12668
rect 24574 11318 24600 11321
rect 24574 11289 24600 11292
rect 24580 11117 24594 11289
rect 24758 11284 24784 11287
rect 24758 11255 24784 11258
rect 24574 11114 24600 11117
rect 24574 11085 24600 11088
rect 24666 10740 24692 10743
rect 24666 10711 24692 10714
rect 24620 10672 24646 10675
rect 24620 10643 24646 10646
rect 24626 10505 24640 10643
rect 24620 10502 24646 10505
rect 24620 10473 24646 10476
rect 24672 10403 24686 10711
rect 24666 10400 24692 10403
rect 24666 10371 24692 10374
rect 24620 9618 24646 9621
rect 24620 9589 24646 9592
rect 24482 8394 24508 8397
rect 24482 8365 24508 8368
rect 24626 8295 24640 9589
rect 24344 8292 24370 8295
rect 24620 8292 24646 8295
rect 24344 8263 24370 8266
rect 24390 8289 24416 8292
rect 24390 8260 24416 8263
rect 24513 8289 24539 8292
rect 24539 8263 24548 8286
rect 24513 8260 24548 8263
rect 24298 8224 24324 8227
rect 24298 8195 24324 8198
rect 24396 8125 24410 8260
rect 24482 8224 24508 8227
rect 24482 8195 24508 8198
rect 24488 8125 24502 8195
rect 24390 8122 24416 8125
rect 24390 8093 24416 8096
rect 24482 8122 24508 8125
rect 24482 8093 24508 8096
rect 23516 8054 23542 8057
rect 23516 8025 23542 8028
rect 23522 7997 23536 8025
rect 23522 7983 23582 7997
rect 23515 7596 23543 7600
rect 23515 7563 23543 7568
rect 23522 7547 23536 7563
rect 23516 7544 23542 7547
rect 23516 7515 23542 7518
rect 23568 7513 23582 7983
rect 24344 7680 24370 7683
rect 24344 7651 24370 7654
rect 23562 7510 23588 7513
rect 23562 7481 23588 7484
rect 23516 7408 23542 7411
rect 23516 7379 23542 7382
rect 23522 7003 23536 7379
rect 23516 7000 23542 7003
rect 23516 6971 23542 6974
rect 23522 6852 23536 6971
rect 23568 6969 23582 7481
rect 24205 7188 24233 7192
rect 24205 7155 24206 7160
rect 24232 7155 24233 7160
rect 24206 7141 24232 7144
rect 23562 6966 23588 6969
rect 23562 6937 23588 6940
rect 23515 6848 23543 6852
rect 23515 6815 23543 6820
rect 23423 6508 23451 6512
rect 23423 6475 23451 6480
rect 23200 6425 23260 6433
rect 23378 6456 23404 6459
rect 23378 6427 23404 6430
rect 23194 6422 23260 6425
rect 23220 6419 23260 6422
rect 23194 6393 23220 6396
rect 22964 6320 22990 6323
rect 22964 6291 22990 6294
rect 22688 5572 22714 5575
rect 22688 5543 22714 5546
rect 22320 5504 22346 5507
rect 22320 5475 22346 5478
rect 22412 5504 22438 5507
rect 22412 5475 22438 5478
rect 22274 5402 22300 5405
rect 22274 5373 22300 5376
rect 22136 5130 22162 5133
rect 22136 5101 22162 5104
rect 21354 4999 21380 5002
rect 21445 5012 21473 5016
rect 21124 4824 21150 4827
rect 21124 4795 21150 4798
rect 21078 4790 21104 4793
rect 21078 4761 21104 4764
rect 21130 4453 21144 4795
rect 21360 4793 21374 4999
rect 21445 4979 21446 4984
rect 21472 4979 21473 4984
rect 21446 4965 21472 4968
rect 22418 4827 22432 5475
rect 23384 5371 23398 6427
rect 23568 6425 23582 6937
rect 24114 6864 24140 6867
rect 24114 6835 24140 6838
rect 23976 6694 24002 6697
rect 23976 6665 24002 6668
rect 23562 6422 23588 6425
rect 23562 6393 23588 6396
rect 23982 6217 23996 6665
rect 24120 6663 24134 6835
rect 24114 6660 24140 6663
rect 24114 6631 24140 6634
rect 24212 6629 24226 7141
rect 24206 6626 24232 6629
rect 24206 6597 24232 6600
rect 24350 6493 24364 7651
rect 24482 7578 24508 7581
rect 24534 7572 24548 8260
rect 24619 8276 24620 8280
rect 24646 8276 24647 8280
rect 24619 8243 24647 8248
rect 24508 7558 24548 7572
rect 24482 7549 24508 7552
rect 24672 7411 24686 10371
rect 24712 8054 24738 8057
rect 24712 8025 24738 8028
rect 24666 7408 24692 7411
rect 24666 7379 24692 7382
rect 24718 6901 24732 8025
rect 24764 7989 24778 11255
rect 24810 10743 24824 12663
rect 25546 12417 25560 12819
rect 25586 12678 25612 12681
rect 25586 12649 25612 12652
rect 25592 12443 25606 12649
rect 25408 12409 25560 12417
rect 25586 12440 25612 12443
rect 25586 12411 25612 12414
rect 25402 12406 25560 12409
rect 25428 12403 25560 12406
rect 25402 12377 25428 12380
rect 25408 12205 25422 12377
rect 25402 12202 25428 12205
rect 25402 12173 25428 12176
rect 25408 11865 25422 12173
rect 25494 12066 25520 12069
rect 25494 12037 25520 12040
rect 25402 11862 25428 11865
rect 25402 11833 25428 11836
rect 25500 11006 25514 12037
rect 25592 11047 25606 12411
rect 25638 12409 25652 12921
rect 25632 12406 25658 12409
rect 25632 12377 25658 12380
rect 25638 12103 25652 12377
rect 25632 12100 25658 12103
rect 25632 12071 25658 12074
rect 25638 11899 25652 12071
rect 25632 11896 25658 11899
rect 25632 11867 25658 11870
rect 25868 11047 25882 12955
rect 26006 12851 26020 13465
rect 26144 12953 26158 13465
rect 26138 12950 26164 12953
rect 26138 12921 26164 12924
rect 26000 12848 26026 12851
rect 26000 12819 26026 12822
rect 26236 12632 26250 13627
rect 26328 13573 26342 15539
rect 26466 14619 26480 17851
rect 26920 17608 26946 17611
rect 26920 17579 26946 17582
rect 26736 17540 26762 17543
rect 26736 17511 26762 17514
rect 26742 17203 26756 17511
rect 26782 17234 26808 17237
rect 26782 17205 26808 17208
rect 26736 17200 26762 17203
rect 26736 17171 26762 17174
rect 26742 16999 26756 17171
rect 26736 16996 26762 16999
rect 26736 16967 26762 16970
rect 26690 16656 26716 16659
rect 26742 16633 26756 16967
rect 26788 16965 26802 17205
rect 26782 16962 26808 16965
rect 26782 16933 26808 16936
rect 26716 16630 26756 16633
rect 26690 16627 26756 16630
rect 26696 16619 26756 16627
rect 26742 16115 26756 16619
rect 26736 16112 26762 16115
rect 26736 16083 26762 16086
rect 26742 15945 26756 16083
rect 26736 15942 26762 15945
rect 26736 15913 26762 15916
rect 26506 15840 26532 15843
rect 26506 15811 26532 15814
rect 26512 15605 26526 15811
rect 26506 15602 26532 15605
rect 26506 15573 26532 15576
rect 26742 15401 26756 15913
rect 26782 15874 26808 15877
rect 26782 15845 26808 15848
rect 26736 15398 26762 15401
rect 26736 15369 26762 15372
rect 26788 15367 26802 15845
rect 26926 15673 26940 17579
rect 27064 17339 27078 18667
rect 27110 18155 27124 21923
rect 27149 21911 27177 21916
rect 27196 21824 27222 21827
rect 27196 21795 27222 21798
rect 27202 20739 27216 21795
rect 27196 20736 27222 20739
rect 27196 20707 27222 20710
rect 27104 18152 27130 18155
rect 27104 18123 27130 18126
rect 27110 17815 27124 18123
rect 27104 17812 27130 17815
rect 27104 17783 27130 17786
rect 27104 17744 27130 17747
rect 27104 17715 27130 17718
rect 27058 17336 27084 17339
rect 27058 17307 27084 17310
rect 26966 17098 26992 17101
rect 26966 17069 26992 17072
rect 26972 16965 26986 17069
rect 26966 16962 26992 16965
rect 26966 16933 26992 16936
rect 27012 15874 27038 15877
rect 27012 15845 27038 15848
rect 26920 15670 26946 15673
rect 26920 15641 26946 15644
rect 26782 15364 26808 15367
rect 26782 15335 26808 15338
rect 26966 15330 26992 15333
rect 26966 15301 26992 15304
rect 26972 15216 26986 15301
rect 26965 15212 26993 15216
rect 26965 15179 26993 15184
rect 26460 14616 26486 14619
rect 26460 14587 26486 14590
rect 26828 14208 26854 14211
rect 26828 14179 26854 14182
rect 26834 13735 26848 14179
rect 26828 13732 26854 13735
rect 26828 13703 26854 13706
rect 26282 13559 26342 13573
rect 26282 12681 26296 13559
rect 27018 13497 27032 15845
rect 27064 13837 27078 17307
rect 27110 17305 27124 17715
rect 27104 17302 27130 17305
rect 27104 17273 27130 17276
rect 27202 16293 27216 20707
rect 27334 20226 27360 20229
rect 27334 20197 27360 20200
rect 27340 19821 27354 20197
rect 27334 19818 27360 19821
rect 27334 19789 27360 19792
rect 27242 19104 27268 19107
rect 27242 19075 27268 19078
rect 27288 19104 27314 19107
rect 27288 19075 27314 19078
rect 27248 17645 27262 19075
rect 27294 18733 27308 19075
rect 27288 18730 27314 18733
rect 27288 18701 27314 18704
rect 27242 17642 27268 17645
rect 27242 17613 27268 17616
rect 27340 17373 27354 19789
rect 27386 19209 27400 21965
rect 28030 21895 28044 22067
rect 28024 21892 28050 21895
rect 28070 21892 28096 21895
rect 28024 21863 28050 21866
rect 28069 21876 28070 21880
rect 28162 21892 28188 21895
rect 28096 21876 28097 21880
rect 28162 21863 28188 21866
rect 28069 21843 28097 21848
rect 28168 21725 28182 21863
rect 28162 21722 28188 21725
rect 28162 21693 28188 21696
rect 28214 21657 28228 22169
rect 28208 21654 28234 21657
rect 28208 21625 28234 21628
rect 28214 20909 28228 21625
rect 28070 20906 28096 20909
rect 28070 20877 28096 20880
rect 28208 20906 28234 20909
rect 28208 20877 28234 20880
rect 28076 20535 28090 20877
rect 28260 20807 28274 22747
rect 28346 22742 28372 22745
rect 28346 22713 28372 22716
rect 28352 22192 28366 22713
rect 29726 22640 29752 22643
rect 29726 22611 29752 22614
rect 28530 22232 28556 22235
rect 28530 22203 28556 22206
rect 28392 22198 28418 22201
rect 28352 22178 28392 22192
rect 28392 22169 28418 22172
rect 28345 21944 28373 21948
rect 28345 21911 28373 21916
rect 28352 21895 28366 21911
rect 28346 21892 28372 21895
rect 28346 21863 28372 21866
rect 28398 21665 28412 22169
rect 28352 21657 28412 21665
rect 28438 21688 28464 21691
rect 28438 21659 28464 21662
rect 28346 21654 28412 21657
rect 28372 21651 28412 21654
rect 28346 21625 28372 21628
rect 28116 20804 28142 20807
rect 28116 20775 28142 20778
rect 28254 20804 28280 20807
rect 28254 20775 28280 20778
rect 28122 20603 28136 20775
rect 28116 20600 28142 20603
rect 28116 20571 28142 20574
rect 28070 20532 28096 20535
rect 28070 20503 28096 20506
rect 28076 20305 28090 20503
rect 28030 20291 28090 20305
rect 28030 20263 28044 20291
rect 28122 20263 28136 20571
rect 28254 20362 28280 20365
rect 28254 20333 28280 20336
rect 28024 20260 28050 20263
rect 28024 20231 28050 20234
rect 28116 20260 28142 20263
rect 28116 20231 28142 20234
rect 27794 20226 27820 20229
rect 27794 20197 27820 20200
rect 27800 19651 27814 20197
rect 27794 19648 27820 19651
rect 27794 19619 27820 19622
rect 27380 19206 27406 19209
rect 27380 19177 27406 19180
rect 28030 18937 28044 20231
rect 28260 20229 28274 20333
rect 28300 20260 28326 20263
rect 28300 20231 28326 20234
rect 28254 20226 28280 20229
rect 28254 20197 28280 20200
rect 28024 18934 28050 18937
rect 27984 18914 28024 18928
rect 27984 18869 27998 18914
rect 28024 18905 28050 18908
rect 28306 18928 28320 20231
rect 28352 19013 28366 21625
rect 28444 20365 28458 21659
rect 28536 20707 28550 22203
rect 29542 22096 29568 22099
rect 29542 22067 29568 22070
rect 29548 21657 29562 22067
rect 29732 21691 29746 22611
rect 29726 21688 29752 21691
rect 29726 21659 29752 21662
rect 29358 21654 29384 21657
rect 29358 21625 29384 21628
rect 29542 21654 29568 21657
rect 29542 21625 29568 21628
rect 29818 21654 29844 21657
rect 29818 21625 29844 21628
rect 29312 21552 29338 21555
rect 29312 21523 29338 21526
rect 28536 20693 28596 20707
rect 28536 20569 28550 20693
rect 28530 20566 28556 20569
rect 28530 20537 28556 20540
rect 28438 20362 28464 20365
rect 28438 20333 28464 20336
rect 28352 18999 28412 19013
rect 28346 18934 28372 18937
rect 28306 18914 28346 18928
rect 27978 18866 28004 18869
rect 27978 18837 28004 18840
rect 27380 18832 27406 18835
rect 27380 18803 27406 18806
rect 27386 18597 27400 18803
rect 27984 18665 27998 18837
rect 27978 18662 28004 18665
rect 27978 18633 28004 18636
rect 27564 18628 27590 18631
rect 27564 18599 27590 18602
rect 27380 18594 27406 18597
rect 27380 18565 27406 18568
rect 27518 18594 27544 18597
rect 27518 18565 27544 18568
rect 27524 18461 27538 18565
rect 27518 18458 27544 18461
rect 27518 18429 27544 18432
rect 27570 18393 27584 18599
rect 27564 18390 27590 18393
rect 27564 18361 27590 18364
rect 27984 18359 27998 18633
rect 28306 18631 28320 18914
rect 28346 18905 28372 18908
rect 28300 18628 28326 18631
rect 28326 18602 28366 18605
rect 28300 18599 28366 18602
rect 28254 18594 28280 18597
rect 28306 18591 28366 18599
rect 28254 18565 28280 18568
rect 28260 18537 28274 18565
rect 28260 18523 28320 18537
rect 27978 18356 28004 18359
rect 27978 18327 28004 18330
rect 27426 17812 27452 17815
rect 27426 17783 27452 17786
rect 27334 17370 27360 17373
rect 27334 17341 27360 17344
rect 27432 17305 27446 17783
rect 27984 17543 27998 18327
rect 28306 18189 28320 18523
rect 28352 18427 28366 18591
rect 28346 18424 28372 18427
rect 28346 18395 28372 18398
rect 28300 18186 28326 18189
rect 28300 18157 28326 18160
rect 27978 17540 28004 17543
rect 27978 17511 28004 17514
rect 27242 17302 27268 17305
rect 27242 17273 27268 17276
rect 27426 17302 27452 17305
rect 27426 17273 27452 17276
rect 27248 16829 27262 17273
rect 27242 16826 27268 16829
rect 27242 16797 27268 16800
rect 27202 16279 27354 16293
rect 27196 16112 27222 16115
rect 27196 16083 27222 16086
rect 27202 15673 27216 16083
rect 27288 15840 27314 15843
rect 27288 15811 27314 15814
rect 27294 15673 27308 15811
rect 27340 15673 27354 16279
rect 27104 15670 27130 15673
rect 27104 15641 27130 15644
rect 27196 15670 27222 15673
rect 27196 15641 27222 15644
rect 27288 15670 27314 15673
rect 27288 15641 27314 15644
rect 27340 15670 27375 15673
rect 27340 15644 27349 15670
rect 27340 15641 27375 15644
rect 27110 15571 27124 15641
rect 27340 15613 27354 15641
rect 27156 15599 27354 15613
rect 27104 15568 27130 15571
rect 27104 15539 27130 15542
rect 27104 14004 27130 14007
rect 27104 13975 27130 13978
rect 27058 13834 27084 13837
rect 27058 13805 27084 13808
rect 26322 13494 26348 13497
rect 26322 13465 26348 13468
rect 27012 13494 27038 13497
rect 27012 13465 27038 13468
rect 26276 12678 26302 12681
rect 26276 12649 26302 12652
rect 26229 12628 26257 12632
rect 26229 12595 26257 12600
rect 26184 11896 26210 11899
rect 26184 11867 26210 11870
rect 26190 11748 26204 11867
rect 26183 11744 26211 11748
rect 26183 11711 26211 11716
rect 25592 11033 25652 11047
rect 25868 11033 25974 11047
rect 25500 10992 25606 11006
rect 25592 10811 25606 10992
rect 25586 10808 25612 10811
rect 25586 10779 25612 10782
rect 24804 10740 24830 10743
rect 24804 10711 24830 10714
rect 25356 10740 25382 10743
rect 25592 10728 25606 10779
rect 25356 10711 25382 10714
rect 25585 10724 25613 10728
rect 24896 10672 24922 10675
rect 24896 10643 24922 10646
rect 24902 10471 24916 10643
rect 24896 10468 24922 10471
rect 24896 10439 24922 10442
rect 25362 10233 25376 10711
rect 25585 10691 25613 10696
rect 25638 10309 25652 11033
rect 25678 10774 25704 10777
rect 25678 10745 25704 10748
rect 25684 10675 25698 10745
rect 25678 10672 25704 10675
rect 25678 10643 25704 10646
rect 25592 10295 25652 10309
rect 25592 10267 25606 10295
rect 25586 10264 25612 10267
rect 25586 10235 25612 10238
rect 25356 10230 25382 10233
rect 25356 10201 25382 10204
rect 25362 9723 25376 10201
rect 25356 9720 25382 9723
rect 25356 9691 25382 9694
rect 25356 9652 25382 9655
rect 25356 9623 25382 9626
rect 25264 9414 25290 9417
rect 25264 9385 25290 9388
rect 24804 8122 24830 8125
rect 24804 8093 24830 8096
rect 24758 7986 24784 7989
rect 24758 7957 24784 7960
rect 24810 7819 24824 8093
rect 25270 8057 25284 9385
rect 25362 9349 25376 9623
rect 25356 9346 25382 9349
rect 25356 9317 25382 9320
rect 25402 9346 25428 9349
rect 25402 9317 25428 9320
rect 25362 9300 25376 9317
rect 25355 9296 25383 9300
rect 25355 9263 25383 9268
rect 25408 9213 25422 9317
rect 25402 9210 25428 9213
rect 25402 9181 25428 9184
rect 25592 8771 25606 10235
rect 25684 10233 25698 10643
rect 25678 10230 25704 10233
rect 25678 10201 25704 10204
rect 25632 9686 25658 9689
rect 25632 9657 25658 9660
rect 25638 9111 25652 9657
rect 25684 9179 25698 10201
rect 25862 9584 25888 9587
rect 25862 9555 25888 9558
rect 25868 9232 25882 9555
rect 25861 9228 25889 9232
rect 25861 9195 25889 9200
rect 25868 9179 25882 9195
rect 25678 9176 25704 9179
rect 25862 9176 25888 9179
rect 25678 9147 25704 9150
rect 25723 9160 25751 9164
rect 25632 9108 25658 9111
rect 25632 9079 25658 9082
rect 25684 8805 25698 9147
rect 25862 9147 25888 9150
rect 25723 9127 25751 9132
rect 25678 8802 25704 8805
rect 25678 8773 25704 8776
rect 25586 8768 25612 8771
rect 25586 8739 25612 8742
rect 25684 8601 25698 8773
rect 25730 8635 25744 9127
rect 25816 9040 25842 9043
rect 25816 9011 25842 9014
rect 25724 8632 25750 8635
rect 25724 8603 25750 8606
rect 25678 8598 25704 8601
rect 25678 8569 25704 8572
rect 25822 8567 25836 9011
rect 25816 8564 25842 8567
rect 25816 8535 25842 8538
rect 25264 8054 25290 8057
rect 25264 8025 25290 8028
rect 24804 7816 24830 7819
rect 24804 7787 24830 7790
rect 25822 7479 25836 8535
rect 25862 7544 25888 7547
rect 25862 7515 25888 7518
rect 25816 7476 25842 7479
rect 25816 7447 25842 7450
rect 25822 7309 25836 7447
rect 25678 7306 25704 7309
rect 25678 7277 25704 7280
rect 25816 7306 25842 7309
rect 25816 7277 25842 7280
rect 24896 7136 24922 7139
rect 24896 7107 24922 7110
rect 24902 7056 24916 7107
rect 24895 7052 24923 7056
rect 24895 7019 24923 7024
rect 24902 6969 24916 7019
rect 24758 6966 24784 6969
rect 24758 6937 24784 6940
rect 24850 6966 24876 6969
rect 24850 6937 24876 6940
rect 24896 6966 24922 6969
rect 24896 6937 24922 6940
rect 24712 6898 24738 6901
rect 24712 6869 24738 6872
rect 24574 6864 24600 6867
rect 24574 6835 24600 6838
rect 24344 6490 24370 6493
rect 24344 6461 24370 6464
rect 24580 6459 24594 6835
rect 24764 6493 24778 6937
rect 24856 6765 24870 6937
rect 25684 6935 25698 7277
rect 25678 6932 25704 6935
rect 25678 6903 25704 6906
rect 24850 6762 24876 6765
rect 24850 6733 24876 6736
rect 24758 6490 24784 6493
rect 24758 6461 24784 6464
rect 24574 6456 24600 6459
rect 24574 6427 24600 6430
rect 25448 6456 25474 6459
rect 25448 6427 25474 6430
rect 23844 6203 23996 6217
rect 23378 5368 23404 5371
rect 23378 5339 23404 5342
rect 23384 5235 23398 5339
rect 23844 5337 23858 6203
rect 24206 5878 24232 5881
rect 24206 5849 24232 5852
rect 24212 5337 24226 5849
rect 25402 5640 25428 5643
rect 25402 5611 25428 5614
rect 25356 5572 25382 5575
rect 25356 5543 25382 5546
rect 25362 5405 25376 5543
rect 25356 5402 25382 5405
rect 25356 5373 25382 5376
rect 25408 5337 25422 5611
rect 25454 5405 25468 6427
rect 25678 5538 25704 5541
rect 25678 5509 25704 5512
rect 25448 5402 25474 5405
rect 25448 5373 25474 5376
rect 25684 5337 25698 5509
rect 23838 5334 23864 5337
rect 23838 5305 23864 5308
rect 24206 5334 24232 5337
rect 25356 5334 25382 5337
rect 24232 5314 24272 5328
rect 24206 5305 24232 5308
rect 23378 5232 23404 5235
rect 23378 5203 23404 5206
rect 23844 5065 23858 5305
rect 23838 5062 23864 5065
rect 23838 5033 23864 5036
rect 22412 4824 22438 4827
rect 22412 4795 22438 4798
rect 21354 4790 21380 4793
rect 21354 4761 21380 4764
rect 23844 4521 23858 5033
rect 24258 5031 24272 5314
rect 25356 5305 25382 5308
rect 25402 5334 25428 5337
rect 25402 5305 25428 5308
rect 25678 5334 25704 5337
rect 25678 5305 25704 5308
rect 25362 5133 25376 5305
rect 25632 5266 25658 5269
rect 25632 5237 25658 5240
rect 25356 5130 25382 5133
rect 25356 5101 25382 5104
rect 24252 5028 24278 5031
rect 24205 5012 24233 5016
rect 24252 4999 24278 5002
rect 24205 4979 24206 4984
rect 24232 4979 24233 4984
rect 24206 4965 24232 4968
rect 24258 4529 24272 4999
rect 25638 4589 25652 5237
rect 25868 5016 25882 7515
rect 25960 7003 25974 11033
rect 26236 10743 26250 12595
rect 26230 10740 26256 10743
rect 26230 10711 26256 10714
rect 26276 10672 26302 10675
rect 26276 10643 26302 10646
rect 26282 10505 26296 10643
rect 26276 10502 26302 10505
rect 26276 10473 26302 10476
rect 26046 10468 26072 10471
rect 26230 10468 26256 10471
rect 26046 10439 26072 10442
rect 26229 10452 26230 10456
rect 26256 10452 26257 10456
rect 26052 10301 26066 10439
rect 26229 10419 26257 10424
rect 26046 10298 26072 10301
rect 26046 10269 26072 10272
rect 26328 7589 26342 13465
rect 26690 12406 26716 12409
rect 26690 12377 26716 12380
rect 26782 12406 26808 12409
rect 26782 12377 26808 12380
rect 26874 12406 26900 12409
rect 26874 12377 26900 12380
rect 26696 11049 26710 12377
rect 26788 12205 26802 12377
rect 26828 12304 26854 12307
rect 26828 12275 26854 12278
rect 26782 12202 26808 12205
rect 26782 12173 26808 12176
rect 26690 11046 26716 11049
rect 26690 11017 26716 11020
rect 26696 10539 26710 11017
rect 26834 10845 26848 12275
rect 26828 10842 26854 10845
rect 26828 10813 26854 10816
rect 26736 10672 26762 10675
rect 26736 10643 26762 10646
rect 26690 10536 26716 10539
rect 26690 10507 26716 10510
rect 26742 9485 26756 10643
rect 26880 10505 26894 12377
rect 27012 10774 27038 10777
rect 27012 10745 27038 10748
rect 26874 10502 26900 10505
rect 26874 10473 26900 10476
rect 26966 9618 26992 9621
rect 26966 9589 26992 9592
rect 26690 9482 26716 9485
rect 26690 9453 26716 9456
rect 26736 9482 26762 9485
rect 26736 9453 26762 9456
rect 26696 9436 26710 9453
rect 26689 9432 26717 9436
rect 26689 9399 26717 9404
rect 26874 9380 26900 9383
rect 26972 9368 26986 9589
rect 26874 9351 26900 9354
rect 26965 9364 26993 9368
rect 26880 9179 26894 9351
rect 26965 9331 26993 9336
rect 26920 9312 26946 9315
rect 26920 9283 26946 9286
rect 26926 9213 26940 9283
rect 26920 9210 26946 9213
rect 26920 9181 26946 9184
rect 26874 9176 26900 9179
rect 26972 9153 26986 9331
rect 26874 9147 26900 9150
rect 26926 9145 26986 9153
rect 26920 9142 26986 9145
rect 26946 9139 26986 9142
rect 26920 9113 26946 9116
rect 26828 8258 26854 8261
rect 26828 8229 26854 8232
rect 26834 7751 26848 8229
rect 26736 7748 26762 7751
rect 26736 7719 26762 7722
rect 26828 7748 26854 7751
rect 26828 7719 26854 7722
rect 26098 7575 26342 7589
rect 26098 7547 26112 7575
rect 26092 7544 26118 7547
rect 26092 7515 26118 7518
rect 26138 7510 26164 7513
rect 26138 7481 26164 7484
rect 26144 7207 26158 7481
rect 26138 7204 26164 7207
rect 26138 7175 26164 7178
rect 25954 7000 25980 7003
rect 25954 6971 25980 6974
rect 25861 5012 25889 5016
rect 25861 4979 25889 4984
rect 25632 4586 25658 4589
rect 25632 4557 25658 4560
rect 23838 4518 23864 4521
rect 23838 4489 23864 4492
rect 24212 4515 24272 4529
rect 24212 4487 24226 4515
rect 25960 4487 25974 6971
rect 26092 6966 26118 6969
rect 26144 6960 26158 7175
rect 26118 6946 26158 6960
rect 26092 6937 26118 6940
rect 26742 6901 26756 7719
rect 26736 6898 26762 6901
rect 26736 6869 26762 6872
rect 26229 6644 26257 6648
rect 26229 6611 26257 6616
rect 26236 5915 26250 6611
rect 26230 5912 26256 5915
rect 26230 5883 26256 5886
rect 26834 5541 26848 7719
rect 26874 7714 26900 7717
rect 26874 7685 26900 7688
rect 26880 7581 26894 7685
rect 26874 7578 26900 7581
rect 26874 7549 26900 7552
rect 26966 7170 26992 7173
rect 26966 7141 26992 7144
rect 26972 6648 26986 7141
rect 26965 6644 26993 6648
rect 26965 6611 26993 6616
rect 27018 5609 27032 10745
rect 27064 9417 27078 13805
rect 27058 9414 27084 9417
rect 27058 9385 27084 9388
rect 27058 9142 27084 9145
rect 27058 9113 27084 9116
rect 27064 8669 27078 9113
rect 27058 8666 27084 8669
rect 27058 8637 27084 8640
rect 27110 7751 27124 13975
rect 27156 13973 27170 15599
rect 27334 15568 27360 15571
rect 27334 15539 27360 15542
rect 27150 13970 27176 13973
rect 27150 13941 27176 13944
rect 27288 13970 27314 13973
rect 27288 13941 27314 13944
rect 27242 13936 27268 13939
rect 27242 13907 27268 13910
rect 27248 13769 27262 13907
rect 27242 13766 27268 13769
rect 27242 13737 27268 13740
rect 27150 13732 27176 13735
rect 27150 13703 27176 13706
rect 27156 12477 27170 13703
rect 27150 12474 27176 12477
rect 27150 12445 27176 12448
rect 27196 12406 27222 12409
rect 27196 12377 27222 12380
rect 27202 11933 27216 12377
rect 27196 11930 27222 11933
rect 27196 11901 27222 11904
rect 27150 10400 27176 10403
rect 27150 10371 27176 10374
rect 27156 9417 27170 10371
rect 27242 9856 27268 9859
rect 27242 9827 27268 9830
rect 27248 9723 27262 9827
rect 27242 9720 27268 9723
rect 27242 9691 27268 9694
rect 27150 9414 27176 9417
rect 27150 9385 27176 9388
rect 27150 9312 27176 9315
rect 27150 9283 27176 9286
rect 27156 8533 27170 9283
rect 27248 9145 27262 9691
rect 27242 9142 27268 9145
rect 27242 9113 27268 9116
rect 27150 8530 27176 8533
rect 27150 8501 27176 8504
rect 27104 7748 27130 7751
rect 27104 7719 27130 7722
rect 27110 6920 27124 7719
rect 27294 7683 27308 13941
rect 27340 13505 27354 15539
rect 27432 14109 27446 17273
rect 27984 17271 27998 17511
rect 28024 17506 28050 17509
rect 28024 17477 28050 17480
rect 28208 17506 28234 17509
rect 28208 17477 28234 17480
rect 28030 17305 28044 17477
rect 28024 17302 28050 17305
rect 28024 17273 28050 17276
rect 27748 17268 27774 17271
rect 27748 17239 27774 17242
rect 27978 17268 28004 17271
rect 27978 17239 28004 17242
rect 27754 17101 27768 17239
rect 27984 17101 27998 17239
rect 27748 17098 27774 17101
rect 27748 17069 27774 17072
rect 27978 17098 28004 17101
rect 27978 17069 28004 17072
rect 28116 16928 28142 16931
rect 28116 16899 28142 16902
rect 27564 15670 27590 15673
rect 27564 15641 27590 15644
rect 27570 15284 27584 15641
rect 27748 15636 27774 15639
rect 27748 15607 27774 15610
rect 27754 15469 27768 15607
rect 28122 15605 28136 16899
rect 28162 15908 28188 15911
rect 28162 15879 28188 15882
rect 28168 15741 28182 15879
rect 28162 15738 28188 15741
rect 28162 15709 28188 15712
rect 28116 15602 28142 15605
rect 28116 15573 28142 15576
rect 27748 15466 27774 15469
rect 27748 15437 27774 15440
rect 27563 15280 27591 15284
rect 27563 15247 27591 15252
rect 27518 14480 27544 14483
rect 27518 14451 27544 14454
rect 27524 14109 27538 14451
rect 27702 14276 27728 14279
rect 27702 14247 27728 14250
rect 27426 14106 27452 14109
rect 27426 14077 27452 14080
rect 27518 14106 27544 14109
rect 27518 14077 27544 14080
rect 27393 14038 27419 14041
rect 27386 14012 27393 14032
rect 27386 14009 27419 14012
rect 27564 14038 27590 14041
rect 27564 14009 27590 14012
rect 27386 13556 27400 14009
rect 27570 13837 27584 14009
rect 27708 14007 27722 14247
rect 27702 14004 27728 14007
rect 27702 13975 27728 13978
rect 28070 14004 28096 14007
rect 28070 13975 28096 13978
rect 27564 13834 27590 13837
rect 27564 13805 27590 13808
rect 27426 13562 27452 13565
rect 27386 13542 27426 13556
rect 27426 13533 27452 13536
rect 27340 13491 27400 13505
rect 27334 12848 27360 12851
rect 27334 12819 27360 12822
rect 27340 12443 27354 12819
rect 27334 12440 27360 12443
rect 27334 12411 27360 12414
rect 27386 12409 27400 13491
rect 28076 12919 28090 13975
rect 28116 12984 28142 12987
rect 28116 12955 28142 12958
rect 27840 12916 27866 12919
rect 27840 12887 27866 12890
rect 28070 12916 28096 12919
rect 28070 12887 28096 12890
rect 27846 12647 27860 12887
rect 28122 12647 28136 12955
rect 28214 12689 28228 17477
rect 28398 17449 28412 18999
rect 28530 18934 28556 18937
rect 28530 18905 28556 18908
rect 28438 18560 28464 18563
rect 28438 18531 28464 18534
rect 28444 18461 28458 18531
rect 28438 18458 28464 18461
rect 28438 18429 28464 18432
rect 28438 18186 28464 18189
rect 28438 18157 28464 18160
rect 28352 17435 28412 17449
rect 28352 17305 28366 17435
rect 28444 17339 28458 18157
rect 28438 17336 28464 17339
rect 28438 17307 28464 17310
rect 28346 17302 28372 17305
rect 28346 17273 28372 17276
rect 28300 16996 28326 16999
rect 28300 16967 28326 16970
rect 28306 16251 28320 16967
rect 28352 16795 28366 17273
rect 28392 17098 28418 17101
rect 28392 17069 28418 17072
rect 28346 16792 28372 16795
rect 28346 16763 28372 16766
rect 28300 16248 28326 16251
rect 28300 16219 28326 16222
rect 28352 16217 28366 16763
rect 28398 16761 28412 17069
rect 28392 16758 28418 16761
rect 28392 16729 28418 16732
rect 28346 16214 28372 16217
rect 28346 16185 28372 16188
rect 28300 16180 28326 16183
rect 28398 16157 28412 16729
rect 28326 16154 28412 16157
rect 28300 16151 28412 16154
rect 28306 16143 28412 16151
rect 28306 15129 28320 16143
rect 28536 15877 28550 18905
rect 28444 15863 28550 15877
rect 28345 15212 28373 15216
rect 28345 15179 28373 15184
rect 28300 15126 28326 15129
rect 28300 15097 28326 15100
rect 28300 15058 28326 15061
rect 28300 15029 28326 15032
rect 28306 14585 28320 15029
rect 28300 14582 28326 14585
rect 28300 14553 28326 14556
rect 28306 14389 28320 14553
rect 28260 14381 28320 14389
rect 28254 14378 28320 14381
rect 28280 14375 28320 14378
rect 28254 14349 28280 14352
rect 28260 14041 28274 14349
rect 28352 14321 28366 15179
rect 28392 15160 28418 15163
rect 28392 15131 28418 15134
rect 28306 14307 28366 14321
rect 28254 14038 28280 14041
rect 28254 14009 28280 14012
rect 28260 12987 28274 14009
rect 28254 12984 28280 12987
rect 28254 12955 28280 12958
rect 28168 12675 28228 12689
rect 28168 12647 28182 12675
rect 27840 12644 27866 12647
rect 27840 12615 27866 12618
rect 28116 12644 28142 12647
rect 28116 12615 28142 12618
rect 28162 12644 28188 12647
rect 28162 12615 28188 12618
rect 27380 12406 27406 12409
rect 27380 12377 27406 12380
rect 27386 8261 27400 12377
rect 27846 12375 27860 12615
rect 28070 12610 28096 12613
rect 28070 12581 28096 12584
rect 27840 12372 27866 12375
rect 27840 12343 27866 12346
rect 27747 10724 27775 10728
rect 27747 10691 27775 10696
rect 27610 10570 27636 10573
rect 27610 10541 27636 10544
rect 27518 10468 27544 10471
rect 27616 10445 27630 10541
rect 27518 10439 27544 10442
rect 27524 10377 27538 10439
rect 27570 10437 27630 10445
rect 27754 10437 27768 10691
rect 27564 10434 27630 10437
rect 27590 10431 27630 10434
rect 27748 10434 27774 10437
rect 27564 10405 27590 10408
rect 27748 10405 27774 10408
rect 27524 10363 27630 10377
rect 27616 10233 27630 10363
rect 27610 10230 27636 10233
rect 27610 10201 27636 10204
rect 27978 10230 28004 10233
rect 27978 10201 28004 10204
rect 27984 9417 27998 10201
rect 28023 9432 28051 9436
rect 27978 9414 28004 9417
rect 28023 9399 28051 9404
rect 27978 9385 28004 9388
rect 27984 9145 27998 9385
rect 28030 9349 28044 9399
rect 28024 9346 28050 9349
rect 28024 9317 28050 9320
rect 28030 9179 28044 9317
rect 28076 9232 28090 12581
rect 28122 12443 28136 12615
rect 28306 12579 28320 14307
rect 28346 14276 28372 14279
rect 28346 14247 28372 14250
rect 28300 12576 28326 12579
rect 28300 12547 28326 12550
rect 28116 12440 28142 12443
rect 28116 12411 28142 12414
rect 28116 12372 28142 12375
rect 28116 12343 28142 12346
rect 28122 11287 28136 12343
rect 28207 11744 28235 11748
rect 28207 11711 28235 11716
rect 28116 11284 28142 11287
rect 28116 11255 28142 11258
rect 28122 10233 28136 11255
rect 28116 10230 28142 10233
rect 28116 10201 28142 10204
rect 28214 9349 28228 11711
rect 28306 9655 28320 12547
rect 28352 11355 28366 14247
rect 28398 13981 28412 15131
rect 28444 14279 28458 15863
rect 28582 15163 28596 20693
rect 29266 20532 29292 20535
rect 29266 20503 29292 20506
rect 29272 19923 29286 20503
rect 29266 19920 29292 19923
rect 29266 19891 29292 19894
rect 28622 19138 28648 19141
rect 28622 19109 28648 19112
rect 28628 18427 28642 19109
rect 28622 18424 28648 18427
rect 28622 18395 28648 18398
rect 28628 17245 28642 18395
rect 28628 17231 28688 17245
rect 28622 17200 28648 17203
rect 28622 17171 28648 17174
rect 28628 17033 28642 17171
rect 28622 17030 28648 17033
rect 28622 17001 28648 17004
rect 28674 16795 28688 17231
rect 28990 16962 29016 16965
rect 28990 16933 29016 16936
rect 28668 16792 28694 16795
rect 28668 16763 28694 16766
rect 28996 15911 29010 16933
rect 29318 15945 29332 21523
rect 29364 20569 29378 21625
rect 29772 21586 29798 21589
rect 29772 21557 29798 21560
rect 29588 20736 29614 20739
rect 29588 20707 29614 20710
rect 29594 20637 29608 20707
rect 29588 20634 29614 20637
rect 29588 20605 29614 20608
rect 29358 20566 29384 20569
rect 29358 20537 29384 20540
rect 29542 20566 29568 20569
rect 29542 20537 29568 20540
rect 29312 15942 29338 15945
rect 29312 15913 29338 15916
rect 28990 15908 29016 15911
rect 28990 15879 29016 15882
rect 28760 15874 28786 15877
rect 28760 15845 28786 15848
rect 28576 15160 28602 15163
rect 28576 15131 28602 15134
rect 28438 14276 28464 14279
rect 28438 14247 28464 14250
rect 28576 14208 28602 14211
rect 28576 14179 28602 14182
rect 28444 14041 28504 14049
rect 28438 14038 28504 14041
rect 28464 14035 28504 14038
rect 28438 14009 28464 14012
rect 28398 13967 28458 13981
rect 28392 12576 28418 12579
rect 28392 12547 28418 12550
rect 28398 12443 28412 12547
rect 28392 12440 28418 12443
rect 28392 12411 28418 12414
rect 28346 11352 28372 11355
rect 28346 11323 28372 11326
rect 28392 11318 28418 11321
rect 28392 11289 28418 11292
rect 28398 10573 28412 11289
rect 28392 10570 28418 10573
rect 28392 10541 28418 10544
rect 28346 10264 28372 10267
rect 28346 10235 28372 10238
rect 28300 9652 28326 9655
rect 28300 9623 28326 9626
rect 28208 9346 28234 9349
rect 28208 9317 28234 9320
rect 28069 9228 28097 9232
rect 28069 9195 28097 9200
rect 28024 9176 28050 9179
rect 28024 9147 28050 9150
rect 27610 9142 27636 9145
rect 27610 9113 27636 9116
rect 27978 9142 28004 9145
rect 27978 9113 28004 9116
rect 27616 8941 27630 9113
rect 27748 9108 27774 9111
rect 27748 9079 27774 9082
rect 27754 8941 27768 9079
rect 27610 8938 27636 8941
rect 27610 8909 27636 8912
rect 27748 8938 27774 8941
rect 27748 8909 27774 8912
rect 27380 8258 27406 8261
rect 27380 8229 27406 8232
rect 27984 8023 27998 9113
rect 28076 9028 28090 9195
rect 28069 9024 28097 9028
rect 28069 8991 28097 8996
rect 28070 8054 28096 8057
rect 28070 8025 28096 8028
rect 27978 8020 28004 8023
rect 27978 7991 28004 7994
rect 27984 7751 27998 7991
rect 28076 7751 28090 8025
rect 27978 7748 28004 7751
rect 27978 7719 28004 7722
rect 28070 7748 28096 7751
rect 28070 7719 28096 7722
rect 27748 7714 27774 7717
rect 27748 7685 27774 7688
rect 27886 7714 27912 7717
rect 27886 7685 27912 7688
rect 27288 7680 27314 7683
rect 27288 7651 27314 7654
rect 27754 7309 27768 7685
rect 27748 7306 27774 7309
rect 27748 7277 27774 7280
rect 27892 7192 27906 7685
rect 27984 7513 27998 7719
rect 27978 7510 28004 7513
rect 27978 7481 28004 7484
rect 27984 7275 27998 7481
rect 27978 7272 28004 7275
rect 27978 7243 28004 7246
rect 27885 7188 27913 7192
rect 27885 7155 27913 7160
rect 27103 6916 27131 6920
rect 27103 6883 27131 6888
rect 27012 5606 27038 5609
rect 27012 5577 27038 5580
rect 27110 5575 27124 6883
rect 27984 6697 27998 7243
rect 28214 6716 28228 9317
rect 28299 9228 28327 9232
rect 28299 9195 28327 9200
rect 28306 7793 28320 9195
rect 28352 8839 28366 10235
rect 28398 10233 28412 10541
rect 28392 10230 28418 10233
rect 28392 10201 28418 10204
rect 28398 9436 28412 10201
rect 28444 9697 28458 13967
rect 28490 9859 28504 14035
rect 28582 13701 28596 14179
rect 28576 13698 28602 13701
rect 28576 13669 28602 13672
rect 28714 13698 28740 13701
rect 28714 13669 28740 13672
rect 28530 12950 28556 12953
rect 28530 12921 28556 12924
rect 28536 11047 28550 12921
rect 28720 11321 28734 13669
rect 28766 13259 28780 15845
rect 29364 14585 29378 20537
rect 29548 20365 29562 20537
rect 29778 20535 29792 21557
rect 29824 21453 29838 21625
rect 29818 21450 29844 21453
rect 29818 21421 29844 21424
rect 29824 20569 29838 21421
rect 29818 20566 29844 20569
rect 29818 20537 29844 20540
rect 29772 20532 29798 20535
rect 29772 20503 29798 20506
rect 29542 20362 29568 20365
rect 29542 20333 29568 20336
rect 29542 19172 29568 19175
rect 29542 19143 29568 19146
rect 29548 18903 29562 19143
rect 29588 18934 29614 18937
rect 29588 18905 29614 18908
rect 29634 18934 29660 18937
rect 29634 18905 29660 18908
rect 29680 18934 29706 18937
rect 29680 18905 29706 18908
rect 29542 18900 29568 18903
rect 29542 18871 29568 18874
rect 29594 17781 29608 18905
rect 29640 18461 29654 18905
rect 29634 18458 29660 18461
rect 29634 18429 29660 18432
rect 29588 17778 29614 17781
rect 29588 17749 29614 17752
rect 29588 17540 29614 17543
rect 29588 17511 29614 17514
rect 29496 17472 29522 17475
rect 29496 17443 29522 17446
rect 29502 17339 29516 17443
rect 29496 17336 29522 17339
rect 29496 17307 29522 17310
rect 29404 17302 29430 17305
rect 29404 17273 29430 17276
rect 29358 14582 29384 14585
rect 29358 14553 29384 14556
rect 28990 13936 29016 13939
rect 28990 13907 29016 13910
rect 28898 13732 28924 13735
rect 28898 13703 28924 13706
rect 28760 13256 28786 13259
rect 28760 13227 28786 13230
rect 28668 11318 28694 11321
rect 28668 11289 28694 11292
rect 28714 11318 28740 11321
rect 28714 11289 28740 11292
rect 28852 11318 28878 11321
rect 28852 11289 28878 11292
rect 28536 11033 28596 11047
rect 28484 9856 28510 9859
rect 28484 9827 28510 9830
rect 28444 9683 28504 9697
rect 28438 9652 28464 9655
rect 28438 9623 28464 9626
rect 28391 9432 28419 9436
rect 28391 9399 28419 9404
rect 28444 9145 28458 9623
rect 28438 9142 28464 9145
rect 28438 9113 28464 9116
rect 28346 8836 28372 8839
rect 28346 8807 28372 8810
rect 28444 8745 28458 9113
rect 28352 8731 28458 8745
rect 28352 8091 28366 8731
rect 28392 8598 28418 8601
rect 28392 8569 28418 8572
rect 28346 8088 28372 8091
rect 28346 8059 28372 8062
rect 28352 7853 28366 8059
rect 28398 8057 28412 8569
rect 28392 8054 28418 8057
rect 28392 8025 28418 8028
rect 28346 7850 28372 7853
rect 28346 7821 28372 7824
rect 28306 7779 28366 7793
rect 28352 7547 28366 7779
rect 28346 7544 28372 7547
rect 28346 7515 28372 7518
rect 28398 7513 28412 8025
rect 28392 7510 28418 7513
rect 28392 7481 28418 7484
rect 28207 6712 28235 6716
rect 27978 6694 28004 6697
rect 28207 6679 28235 6684
rect 27978 6665 28004 6668
rect 27984 6425 27998 6665
rect 28214 6629 28228 6679
rect 28398 6663 28412 7481
rect 28392 6660 28418 6663
rect 28392 6631 28418 6634
rect 28208 6626 28234 6629
rect 28208 6597 28234 6600
rect 28398 6501 28412 6631
rect 28490 6512 28504 9683
rect 28582 7600 28596 11033
rect 28622 9856 28648 9859
rect 28622 9827 28648 9830
rect 28628 7751 28642 9827
rect 28674 9587 28688 11289
rect 28858 9621 28872 11289
rect 28852 9618 28878 9621
rect 28852 9589 28878 9592
rect 28668 9584 28694 9587
rect 28668 9555 28694 9558
rect 28805 9500 28833 9504
rect 28805 9467 28833 9472
rect 28812 8635 28826 9467
rect 28806 8632 28832 8635
rect 28806 8603 28832 8606
rect 28904 8601 28918 13703
rect 28996 13701 29010 13907
rect 28990 13698 29016 13701
rect 28990 13669 29016 13672
rect 29082 11114 29108 11117
rect 29082 11085 29108 11088
rect 29088 10845 29102 11085
rect 29082 10842 29108 10845
rect 29082 10813 29108 10816
rect 28944 10774 28970 10777
rect 28944 10745 28970 10748
rect 28950 10505 28964 10745
rect 28944 10502 28970 10505
rect 28944 10473 28970 10476
rect 28990 10468 29016 10471
rect 28990 10439 29016 10442
rect 28996 9723 29010 10439
rect 29128 10434 29154 10437
rect 29128 10405 29154 10408
rect 29134 10301 29148 10405
rect 29128 10298 29154 10301
rect 29128 10269 29154 10272
rect 28990 9720 29016 9723
rect 28990 9691 29016 9694
rect 29036 9482 29062 9485
rect 29036 9453 29062 9456
rect 28990 8632 29016 8635
rect 28990 8603 29016 8606
rect 28898 8598 28924 8601
rect 28898 8569 28924 8572
rect 28622 7748 28648 7751
rect 28622 7719 28648 7722
rect 28575 7596 28603 7600
rect 28575 7563 28603 7568
rect 28352 6487 28412 6501
rect 28483 6508 28511 6512
rect 28352 6425 28366 6487
rect 28483 6475 28511 6480
rect 28490 6459 28504 6475
rect 28484 6456 28510 6459
rect 28484 6427 28510 6430
rect 27978 6422 28004 6425
rect 27978 6393 28004 6396
rect 28208 6422 28234 6425
rect 28208 6393 28234 6396
rect 28346 6422 28372 6425
rect 28346 6393 28372 6396
rect 28214 5813 28228 6393
rect 28352 5881 28366 6393
rect 28582 5915 28596 7563
rect 28904 7056 28918 8569
rect 28996 7853 29010 8603
rect 29042 7853 29056 9453
rect 29174 9380 29200 9383
rect 29174 9351 29200 9354
rect 29128 8564 29154 8567
rect 29128 8535 29154 8538
rect 29134 8125 29148 8535
rect 29128 8122 29154 8125
rect 29128 8093 29154 8096
rect 29180 8065 29194 9351
rect 29364 8295 29378 14553
rect 29410 12953 29424 17273
rect 29496 17200 29522 17203
rect 29496 17171 29522 17174
rect 29502 16999 29516 17171
rect 29496 16996 29522 16999
rect 29496 16967 29522 16970
rect 29496 16928 29522 16931
rect 29496 16899 29522 16902
rect 29502 16557 29516 16899
rect 29496 16554 29522 16557
rect 29496 16525 29522 16528
rect 29594 16455 29608 17511
rect 29634 16656 29660 16659
rect 29634 16627 29660 16630
rect 29640 16455 29654 16627
rect 29686 16455 29700 18905
rect 29772 18390 29798 18393
rect 29772 18361 29798 18364
rect 29778 17305 29792 18361
rect 29772 17302 29798 17305
rect 29772 17273 29798 17276
rect 29588 16452 29614 16455
rect 29588 16423 29614 16426
rect 29634 16452 29660 16455
rect 29634 16423 29660 16426
rect 29680 16452 29706 16455
rect 29680 16423 29706 16426
rect 29818 16452 29844 16455
rect 29818 16423 29844 16426
rect 29496 16418 29522 16421
rect 29496 16389 29522 16392
rect 29502 16285 29516 16389
rect 29496 16282 29522 16285
rect 29496 16253 29522 16256
rect 29725 15280 29753 15284
rect 29725 15247 29753 15252
rect 29450 15024 29476 15027
rect 29450 14995 29476 14998
rect 29456 14585 29470 14995
rect 29450 14582 29476 14585
rect 29450 14553 29476 14556
rect 29588 14480 29614 14483
rect 29588 14451 29614 14454
rect 29594 13735 29608 14451
rect 29496 13732 29522 13735
rect 29496 13703 29522 13706
rect 29588 13732 29614 13735
rect 29588 13703 29614 13706
rect 29502 13021 29516 13703
rect 29542 13664 29568 13667
rect 29542 13635 29568 13638
rect 29548 13293 29562 13635
rect 29542 13290 29568 13293
rect 29542 13261 29568 13264
rect 29496 13018 29522 13021
rect 29496 12989 29522 12992
rect 29732 12953 29746 15247
rect 29824 12953 29838 16423
rect 31749 15280 31777 15284
rect 31749 15247 31777 15252
rect 31756 15061 31770 15247
rect 31750 15058 31776 15061
rect 31750 15029 31776 15032
rect 29404 12950 29430 12953
rect 29404 12921 29430 12924
rect 29542 12950 29568 12953
rect 29542 12921 29568 12924
rect 29634 12950 29660 12953
rect 29634 12921 29660 12924
rect 29709 12950 29746 12953
rect 29735 12924 29746 12950
rect 29709 12921 29746 12924
rect 29818 12950 29844 12953
rect 29818 12921 29844 12924
rect 29410 9655 29424 12921
rect 29548 12749 29562 12921
rect 29640 12893 29654 12921
rect 29640 12879 29700 12893
rect 29542 12746 29568 12749
rect 29542 12717 29568 12720
rect 29686 12409 29700 12879
rect 29680 12406 29706 12409
rect 29680 12377 29706 12380
rect 29588 12304 29614 12307
rect 29588 12275 29614 12278
rect 29450 11216 29476 11219
rect 29450 11187 29476 11190
rect 29456 10777 29470 11187
rect 29496 10808 29522 10811
rect 29496 10779 29522 10782
rect 29450 10774 29476 10777
rect 29450 10745 29476 10748
rect 29404 9652 29430 9655
rect 29404 9623 29430 9626
rect 29358 8292 29384 8295
rect 29358 8263 29384 8266
rect 29134 8051 29194 8065
rect 28990 7850 29016 7853
rect 28990 7821 29016 7824
rect 29036 7850 29062 7853
rect 29036 7821 29062 7824
rect 28897 7052 28925 7056
rect 28897 7019 28925 7024
rect 29134 7003 29148 8051
rect 29312 7748 29338 7751
rect 29312 7719 29338 7722
rect 29128 7000 29154 7003
rect 29127 6984 29128 6988
rect 29154 6984 29155 6988
rect 29036 6966 29062 6969
rect 29127 6951 29155 6956
rect 29174 6966 29200 6969
rect 29036 6937 29062 6940
rect 29174 6937 29200 6940
rect 29042 6765 29056 6937
rect 29036 6762 29062 6765
rect 29036 6733 29062 6736
rect 29180 6391 29194 6937
rect 29318 6901 29332 7719
rect 29364 6969 29378 8263
rect 29410 7717 29424 9623
rect 29502 9485 29516 10779
rect 29496 9482 29522 9485
rect 29496 9453 29522 9456
rect 29594 9383 29608 12275
rect 29732 9667 29746 12921
rect 29686 9653 29746 9667
rect 29686 9504 29700 9653
rect 29679 9500 29707 9504
rect 29679 9467 29707 9472
rect 29686 9383 29700 9467
rect 29588 9380 29614 9383
rect 29588 9351 29614 9354
rect 29680 9380 29706 9383
rect 29680 9351 29706 9354
rect 29634 9346 29660 9349
rect 29634 9317 29660 9320
rect 29640 9213 29654 9317
rect 29634 9210 29660 9213
rect 29634 9181 29660 9184
rect 29725 8276 29753 8280
rect 29824 8269 29838 12921
rect 29753 8255 29838 8269
rect 29725 8243 29753 8248
rect 29732 7751 29746 8243
rect 29542 7748 29568 7751
rect 29542 7719 29568 7722
rect 29726 7748 29752 7751
rect 29726 7719 29752 7722
rect 29404 7714 29430 7717
rect 29404 7685 29430 7688
rect 29548 7581 29562 7719
rect 29680 7714 29706 7717
rect 29680 7685 29706 7688
rect 29542 7578 29568 7581
rect 29542 7549 29568 7552
rect 29358 6966 29384 6969
rect 29358 6937 29384 6940
rect 29312 6898 29338 6901
rect 29312 6869 29338 6872
rect 29174 6388 29200 6391
rect 29174 6359 29200 6362
rect 29686 5949 29700 7685
rect 29680 5946 29706 5949
rect 29680 5917 29706 5920
rect 28576 5912 28602 5915
rect 28576 5883 28602 5886
rect 28346 5878 28372 5881
rect 28346 5849 28372 5852
rect 28208 5810 28234 5813
rect 28208 5781 28234 5784
rect 27288 5776 27314 5779
rect 27288 5747 27314 5750
rect 27294 5575 27308 5747
rect 27104 5572 27130 5575
rect 27104 5543 27130 5546
rect 27288 5572 27314 5575
rect 27288 5543 27314 5546
rect 26828 5538 26854 5541
rect 26828 5509 26854 5512
rect 24206 4484 24232 4487
rect 24206 4455 24232 4458
rect 25954 4484 25980 4487
rect 25954 4455 25980 4458
rect 21124 4450 21150 4453
rect 21124 4421 21150 4424
rect 18778 3940 18804 3943
rect 18778 3911 18804 3914
rect 20388 3940 20414 3943
rect 20388 3911 20414 3914
rect 18646 1373 18706 1387
rect 16294 676 16320 679
rect 16294 647 16320 650
rect 16708 676 16734 679
rect 16708 647 16734 650
rect 16300 0 16314 647
rect 18692 0 18706 1373
rect 18784 0 18798 3911
<< via2 >>
rect 3367 24034 3395 24052
rect 3367 24024 3368 24034
rect 3368 24024 3394 24034
rect 3394 24024 3395 24034
rect 3137 16214 3165 16232
rect 3137 16204 3138 16214
rect 3138 16204 3164 16214
rect 3164 16204 3165 16214
rect 4885 24636 4913 24664
rect 5115 24636 5143 24664
rect 4977 22410 4978 22420
rect 4978 22410 5004 22420
rect 5004 22410 5005 22420
rect 4977 22392 5005 22410
rect 4931 19410 4959 19428
rect 4931 19400 4932 19410
rect 4932 19400 4958 19410
rect 4958 19400 4959 19410
rect 4839 18516 4867 18544
rect 5207 24568 5235 24596
rect 5161 22392 5189 22420
rect 5023 18380 5051 18408
rect 4287 16282 4315 16300
rect 4287 16272 4288 16282
rect 4288 16272 4314 16282
rect 4314 16272 4315 16282
rect 4517 16214 4545 16232
rect 4517 16204 4518 16214
rect 4518 16204 4544 16214
rect 4544 16204 4545 16214
rect 4747 16426 4748 16436
rect 4748 16426 4774 16436
rect 4774 16426 4775 16436
rect 4747 16408 4775 16426
rect 4931 16272 4959 16300
rect 4747 13280 4775 13308
rect 4885 14504 4913 14532
rect 3413 12610 3441 12628
rect 3413 12600 3414 12610
rect 3414 12600 3440 12610
rect 3440 12600 3441 12610
rect 5529 19400 5557 19428
rect 5759 20770 5787 20788
rect 5759 20760 5760 20770
rect 5760 20760 5786 20770
rect 5786 20760 5787 20770
rect 5851 20760 5879 20788
rect 5391 11988 5419 12016
rect 6587 28726 6615 28744
rect 6587 28716 6588 28726
rect 6588 28716 6614 28726
rect 6614 28716 6615 28726
rect 6955 23956 6983 23984
rect 6495 22392 6523 22420
rect 6817 21110 6845 21128
rect 6817 21100 6818 21110
rect 6818 21100 6844 21110
rect 6844 21100 6845 21110
rect 7001 19672 7029 19700
rect 5989 16272 6017 16300
rect 6771 16408 6799 16436
rect 6035 14572 6063 14600
rect 6817 14582 6845 14600
rect 6817 14572 6818 14582
rect 6818 14572 6844 14582
rect 6844 14572 6845 14582
rect 7139 15116 7167 15144
rect 7185 13280 7213 13308
rect 6909 12464 6937 12492
rect 6863 11444 6891 11472
rect 7599 15116 7627 15144
rect 8243 24586 8244 24596
rect 8244 24586 8270 24596
rect 8270 24586 8271 24596
rect 8243 24568 8271 24586
rect 8381 24024 8409 24052
rect 8887 23498 8888 23508
rect 8888 23498 8914 23508
rect 8914 23498 8915 23508
rect 8887 23480 8915 23498
rect 8703 19682 8731 19700
rect 8703 19672 8704 19682
rect 8704 19672 8730 19682
rect 8730 19672 8731 19682
rect 9669 23956 9697 23984
rect 9899 21780 9927 21808
rect 9025 16272 9053 16300
rect 7783 14572 7811 14600
rect 7921 14504 7949 14532
rect 9531 18400 9559 18408
rect 9531 18380 9547 18400
rect 9547 18380 9559 18400
rect 10543 24636 10571 24664
rect 10267 22800 10295 22828
rect 10359 21916 10387 21944
rect 10221 20760 10249 20788
rect 10773 18602 10774 18612
rect 10774 18602 10800 18612
rect 10800 18602 10801 18612
rect 10773 18584 10801 18602
rect 11555 22052 11583 22080
rect 11095 21100 11123 21128
rect 11141 20828 11169 20856
rect 11279 20828 11307 20856
rect 11877 21440 11905 21468
rect 11923 20022 11951 20040
rect 11923 20012 11924 20022
rect 11924 20012 11950 20022
rect 11950 20012 11951 20022
rect 11187 19682 11215 19700
rect 11187 19672 11188 19682
rect 11188 19672 11214 19682
rect 11214 19672 11215 19682
rect 10819 18380 10847 18408
rect 8197 13212 8225 13240
rect 8105 13162 8115 13172
rect 8115 13162 8133 13172
rect 7599 12396 7627 12424
rect 8105 13144 8133 13162
rect 7921 12396 7949 12424
rect 8749 13698 8777 13716
rect 8749 13688 8750 13698
rect 8750 13688 8776 13698
rect 8776 13688 8777 13698
rect 8979 13348 9007 13376
rect 7323 11920 7351 11948
rect 9025 12600 9053 12628
rect 12015 24296 12043 24324
rect 12383 21110 12411 21128
rect 12383 21100 12384 21110
rect 12384 21100 12410 21110
rect 12410 21100 12411 21110
rect 12383 20216 12411 20244
rect 12245 16970 12246 16980
rect 12246 16970 12272 16980
rect 12272 16970 12273 16980
rect 12245 16952 12273 16970
rect 11739 16758 11767 16776
rect 11739 16748 11740 16758
rect 11740 16748 11766 16758
rect 11766 16748 11767 16758
rect 11187 16272 11215 16300
rect 9669 12124 9697 12152
rect 9117 11862 9145 11880
rect 9117 11852 9118 11862
rect 9118 11852 9144 11862
rect 9144 11852 9145 11862
rect 8795 11784 8823 11812
rect 9577 11716 9605 11744
rect 8703 11444 8731 11472
rect 10083 13290 10111 13308
rect 10083 13280 10084 13290
rect 10084 13280 10110 13290
rect 10110 13280 10111 13290
rect 9991 11920 10019 11948
rect 12107 15116 12135 15144
rect 10267 13552 10295 13580
rect 10911 13698 10939 13716
rect 10911 13688 10912 13698
rect 10912 13688 10938 13698
rect 10938 13688 10939 13698
rect 11739 13280 11767 13308
rect 11739 13144 11767 13172
rect 10405 12474 10433 12492
rect 10405 12464 10406 12474
rect 10406 12464 10432 12474
rect 10432 12464 10433 12474
rect 12613 19962 12614 19972
rect 12614 19962 12640 19972
rect 12640 19962 12641 19972
rect 12613 19944 12641 19962
rect 12061 13212 12089 13240
rect 12659 18584 12687 18612
rect 12889 21780 12917 21808
rect 12383 14504 12411 14532
rect 11647 12406 11675 12424
rect 11647 12396 11648 12406
rect 11648 12396 11674 12406
rect 11674 12396 11675 12406
rect 12015 12124 12043 12152
rect 11739 11852 11767 11880
rect 11049 11784 11077 11812
rect 11647 11784 11675 11812
rect 11923 11716 11951 11744
rect 12935 21110 12963 21128
rect 12935 21100 12936 21110
rect 12936 21100 12962 21110
rect 12962 21100 12963 21110
rect 13119 19944 13147 19972
rect 12889 17020 12917 17048
rect 13119 18602 13120 18612
rect 13120 18602 13146 18612
rect 13146 18602 13147 18612
rect 13119 18584 13147 18602
rect 13855 24296 13883 24324
rect 13901 23480 13929 23508
rect 13625 18108 13653 18136
rect 13165 16816 13193 16844
rect 14223 28716 14251 28744
rect 14085 20216 14113 20244
rect 13257 14504 13285 14532
rect 13027 11920 13055 11948
rect 14039 13688 14067 13716
rect 14223 20012 14251 20040
rect 14407 20234 14423 20244
rect 14423 20234 14435 20244
rect 14407 20216 14435 20234
rect 14131 13620 14159 13648
rect 13855 12396 13883 12424
rect 13165 12328 13193 12356
rect 14591 18108 14619 18136
rect 15097 22052 15125 22080
rect 14913 18584 14941 18612
rect 14637 16758 14665 16776
rect 14637 16748 14638 16758
rect 14638 16748 14664 16758
rect 14664 16748 14665 16758
rect 14545 16690 14573 16708
rect 14545 16680 14546 16690
rect 14546 16680 14572 16690
rect 14572 16680 14573 16690
rect 14545 15116 14573 15144
rect 14545 13688 14573 13716
rect 14729 13552 14757 13580
rect 14637 13162 14638 13172
rect 14638 13162 14664 13172
rect 14664 13162 14665 13172
rect 14637 13144 14665 13162
rect 15603 22052 15631 22080
rect 15189 21440 15217 21468
rect 15143 16970 15144 16980
rect 15144 16970 15170 16980
rect 15170 16970 15171 16980
rect 15143 16952 15171 16970
rect 14959 13280 14987 13308
rect 14499 12124 14527 12152
rect 14407 11852 14435 11880
rect 14361 11716 14389 11744
rect 7139 7568 7167 7596
rect 5207 5596 5235 5624
rect 8749 7654 8750 7664
rect 8750 7654 8776 7664
rect 8776 7654 8777 7664
rect 8749 7636 8777 7654
rect 8841 7568 8869 7596
rect 5529 632 5557 660
rect 15557 16816 15585 16844
rect 15511 16758 15539 16776
rect 15511 16748 15512 16758
rect 15512 16748 15538 16758
rect 15538 16748 15539 16758
rect 17259 26404 17287 26432
rect 16431 21916 16459 21944
rect 16017 16962 16045 16980
rect 16017 16952 16018 16962
rect 16018 16952 16044 16962
rect 16044 16952 16045 16962
rect 15971 16758 15999 16776
rect 15971 16748 15972 16758
rect 15972 16748 15998 16758
rect 15998 16748 15999 16758
rect 15373 13552 15401 13580
rect 15281 12328 15309 12356
rect 15465 11920 15493 11948
rect 17121 22800 17149 22828
rect 16477 16952 16505 16980
rect 16293 13620 16321 13648
rect 17121 16680 17149 16708
rect 18639 26404 18667 26432
rect 18317 13494 18345 13512
rect 18317 13484 18318 13494
rect 18318 13484 18344 13494
rect 18344 13484 18345 13494
rect 17075 10356 17103 10384
rect 16707 9608 16735 9636
rect 18685 18448 18713 18476
rect 18639 15728 18667 15756
rect 18915 18448 18943 18476
rect 19053 13494 19081 13512
rect 19053 13484 19054 13494
rect 19054 13484 19080 13494
rect 19080 13484 19081 13494
rect 19237 12958 19238 12968
rect 19238 12958 19264 12968
rect 19264 12958 19265 12968
rect 19237 12940 19265 12958
rect 20755 19944 20783 19972
rect 20341 18516 20369 18544
rect 20111 16884 20139 16912
rect 20617 18516 20645 18544
rect 20433 12610 20461 12628
rect 20433 12600 20434 12610
rect 20434 12600 20460 12610
rect 20460 12600 20461 12610
rect 20433 9472 20461 9500
rect 20571 6820 20599 6848
rect 20939 18380 20967 18408
rect 20985 15728 21013 15756
rect 21307 22324 21335 22352
rect 21261 16612 21289 16640
rect 20939 9200 20967 9228
rect 21629 18584 21657 18612
rect 21353 16612 21381 16640
rect 22457 18516 22485 18544
rect 22043 17506 22071 17524
rect 22043 17496 22044 17506
rect 22044 17496 22070 17506
rect 22070 17496 22071 17506
rect 22687 16884 22715 16912
rect 21353 10832 21381 10860
rect 21353 9268 21381 9296
rect 21629 12668 21657 12696
rect 21261 6684 21289 6712
rect 21307 6480 21335 6508
rect 21951 6956 21979 6984
rect 21445 6548 21473 6576
rect 22917 19944 22945 19972
rect 22917 19536 22945 19564
rect 23055 18448 23083 18476
rect 23239 17360 23267 17388
rect 22411 9336 22439 9364
rect 22687 10424 22715 10452
rect 22595 6888 22623 6916
rect 22917 10774 22945 10792
rect 22917 10764 22918 10774
rect 22918 10764 22944 10774
rect 22944 10764 22945 10774
rect 23377 10764 23405 10792
rect 23975 17496 24003 17524
rect 23929 12940 23957 12968
rect 23515 10842 23543 10860
rect 23515 10832 23516 10842
rect 23516 10832 23542 10842
rect 23542 10832 23543 10842
rect 22963 9336 22991 9364
rect 24435 22324 24463 22352
rect 24389 19536 24417 19564
rect 24481 18594 24509 18612
rect 24481 18584 24482 18594
rect 24482 18584 24508 18594
rect 24508 18584 24509 18594
rect 24481 18390 24509 18408
rect 24481 18380 24482 18390
rect 24482 18380 24508 18390
rect 24508 18380 24509 18390
rect 23423 10424 23451 10452
rect 23883 9150 23884 9160
rect 23884 9150 23910 9160
rect 23910 9150 23911 9160
rect 23883 9132 23911 9150
rect 24205 9014 24206 9024
rect 24206 9014 24232 9024
rect 24232 9014 24233 9024
rect 24205 8996 24233 9014
rect 25861 21866 25862 21876
rect 25862 21866 25888 21876
rect 25888 21866 25889 21876
rect 25861 21848 25889 21866
rect 25585 17360 25613 17388
rect 25907 17360 25935 17388
rect 26137 16612 26165 16640
rect 24803 12668 24831 12696
rect 23515 7568 23543 7596
rect 24205 7170 24233 7188
rect 24205 7160 24206 7170
rect 24206 7160 24232 7170
rect 24232 7160 24233 7170
rect 23515 6820 23543 6848
rect 23423 6480 23451 6508
rect 21445 4994 21473 5012
rect 21445 4984 21446 4994
rect 21446 4984 21472 4994
rect 21472 4984 21473 4994
rect 24619 8266 24620 8276
rect 24620 8266 24646 8276
rect 24646 8266 24647 8276
rect 24619 8248 24647 8266
rect 27149 21916 27177 21944
rect 26965 15184 26993 15212
rect 28069 21866 28070 21876
rect 28070 21866 28096 21876
rect 28096 21866 28097 21876
rect 28069 21848 28097 21866
rect 28345 21916 28373 21944
rect 26229 12600 26257 12628
rect 26183 11716 26211 11744
rect 25585 10696 25613 10724
rect 25355 9268 25383 9296
rect 25861 9200 25889 9228
rect 25723 9132 25751 9160
rect 24895 7024 24923 7052
rect 24205 4994 24233 5012
rect 24205 4984 24206 4994
rect 24206 4984 24232 4994
rect 24232 4984 24233 4994
rect 26229 10442 26230 10452
rect 26230 10442 26256 10452
rect 26256 10442 26257 10452
rect 26229 10424 26257 10442
rect 26689 9404 26717 9432
rect 26965 9336 26993 9364
rect 25861 4984 25889 5012
rect 26229 6616 26257 6644
rect 26965 6616 26993 6644
rect 27563 15252 27591 15280
rect 28345 15184 28373 15212
rect 27747 10696 27775 10724
rect 28023 9404 28051 9432
rect 28207 11716 28235 11744
rect 28069 9200 28097 9228
rect 28069 8996 28097 9024
rect 27885 7160 27913 7188
rect 27103 6888 27131 6916
rect 28299 9200 28327 9228
rect 28391 9404 28419 9432
rect 28207 6684 28235 6712
rect 28805 9472 28833 9500
rect 28575 7568 28603 7596
rect 28483 6480 28511 6508
rect 29725 15252 29753 15280
rect 31749 15252 31777 15280
rect 28897 7024 28925 7052
rect 29127 6974 29128 6984
rect 29128 6974 29154 6984
rect 29154 6974 29155 6984
rect 29127 6956 29155 6974
rect 29679 9472 29707 9500
rect 29725 8248 29753 8276
<< metal3 >>
rect 6584 28745 6617 28746
rect 14220 28745 14253 28746
rect 6584 28744 14253 28745
rect 6584 28716 6587 28744
rect 6615 28716 14223 28744
rect 14251 28716 14253 28744
rect 6584 28715 14253 28716
rect 6584 28713 6617 28715
rect 14220 28713 14253 28715
rect 17256 26433 17289 26434
rect 18636 26433 18669 26434
rect 17256 26432 18669 26433
rect 17256 26404 17259 26432
rect 17287 26404 18639 26432
rect 18667 26404 18669 26432
rect 17256 26403 18669 26404
rect 17256 26401 17289 26403
rect 18636 26401 18669 26403
rect 4882 24665 4915 24666
rect 5112 24665 5145 24666
rect 10540 24665 10573 24666
rect 4882 24664 10573 24665
rect 4882 24636 4885 24664
rect 4913 24636 5115 24664
rect 5143 24636 10543 24664
rect 10571 24636 10573 24664
rect 4882 24635 10573 24636
rect 4882 24633 4915 24635
rect 5112 24633 5145 24635
rect 10540 24633 10573 24635
rect 5204 24597 5237 24598
rect 8240 24597 8273 24598
rect 5204 24596 8273 24597
rect 5204 24568 5207 24596
rect 5235 24568 8243 24596
rect 8271 24568 8273 24596
rect 5204 24567 8273 24568
rect 5204 24565 5237 24567
rect 8240 24565 8273 24567
rect 12012 24325 12045 24326
rect 13852 24325 13885 24326
rect 12012 24324 13885 24325
rect 12012 24296 12015 24324
rect 12043 24296 13855 24324
rect 13883 24296 13885 24324
rect 12012 24295 13885 24296
rect 12012 24293 12045 24295
rect 13852 24293 13885 24295
rect 3364 24053 3397 24054
rect 8378 24053 8411 24054
rect 3364 24052 8411 24053
rect 3364 24024 3367 24052
rect 3395 24024 8381 24052
rect 8409 24024 8411 24052
rect 3364 24023 8411 24024
rect 3364 24021 3397 24023
rect 8378 24021 8411 24023
rect 6952 23985 6985 23986
rect 9666 23985 9699 23986
rect 6952 23984 9699 23985
rect 6952 23956 6955 23984
rect 6983 23956 9669 23984
rect 9697 23956 9699 23984
rect 6952 23955 9699 23956
rect 6952 23953 6985 23955
rect 9666 23953 9699 23955
rect 8884 23509 8917 23510
rect 13898 23509 13931 23510
rect 8884 23508 13931 23509
rect 8884 23480 8887 23508
rect 8915 23480 13901 23508
rect 13929 23480 13931 23508
rect 8884 23479 13931 23480
rect 8884 23477 8917 23479
rect 13898 23477 13931 23479
rect 10264 22829 10297 22830
rect 17118 22829 17151 22830
rect 10264 22828 17151 22829
rect 10264 22800 10267 22828
rect 10295 22800 17121 22828
rect 17149 22800 17151 22828
rect 10264 22799 17151 22800
rect 10264 22797 10297 22799
rect 17118 22797 17151 22799
rect 4974 22421 5007 22422
rect 5158 22421 5191 22422
rect 6492 22421 6525 22422
rect 4974 22420 6525 22421
rect 4974 22392 4977 22420
rect 5005 22392 5161 22420
rect 5189 22392 6495 22420
rect 6523 22392 6525 22420
rect 4974 22391 6525 22392
rect 4974 22389 5007 22391
rect 5158 22389 5191 22391
rect 6492 22389 6525 22391
rect 21304 22353 21337 22354
rect 24432 22353 24465 22354
rect 21304 22352 24465 22353
rect 21304 22324 21307 22352
rect 21335 22324 24435 22352
rect 24463 22324 24465 22352
rect 21304 22323 24465 22324
rect 21304 22321 21337 22323
rect 24432 22321 24465 22323
rect 11552 22081 11585 22082
rect 15094 22081 15127 22082
rect 15600 22081 15633 22082
rect 11552 22080 15633 22081
rect 11552 22052 11555 22080
rect 11583 22052 15097 22080
rect 15125 22052 15603 22080
rect 15631 22052 15633 22080
rect 11552 22051 15633 22052
rect 11552 22049 11585 22051
rect 15094 22049 15127 22051
rect 15600 22049 15633 22051
rect 10356 21945 10389 21946
rect 16428 21945 16461 21946
rect 10356 21944 16461 21945
rect 10356 21916 10359 21944
rect 10387 21916 16431 21944
rect 16459 21916 16461 21944
rect 10356 21915 16461 21916
rect 10356 21913 10389 21915
rect 16428 21913 16461 21915
rect 27146 21945 27179 21946
rect 28342 21945 28375 21946
rect 27146 21944 28375 21945
rect 27146 21916 27149 21944
rect 27177 21916 28345 21944
rect 28373 21916 28375 21944
rect 27146 21915 28375 21916
rect 27146 21913 27179 21915
rect 28342 21913 28375 21915
rect 25858 21877 25891 21878
rect 28066 21877 28099 21878
rect 25858 21876 28099 21877
rect 25858 21848 25861 21876
rect 25889 21848 28069 21876
rect 28097 21848 28099 21876
rect 25858 21847 28099 21848
rect 25858 21845 25891 21847
rect 28066 21845 28099 21847
rect 9896 21809 9929 21810
rect 12886 21809 12919 21810
rect 9896 21808 12919 21809
rect 9896 21780 9899 21808
rect 9927 21780 12889 21808
rect 12917 21780 12919 21808
rect 9896 21779 12919 21780
rect 9896 21777 9929 21779
rect 12886 21777 12919 21779
rect 11874 21469 11907 21470
rect 15186 21469 15219 21470
rect 11874 21468 15219 21469
rect 11874 21440 11877 21468
rect 11905 21440 15189 21468
rect 15217 21440 15219 21468
rect 11874 21439 15219 21440
rect 11874 21437 11907 21439
rect 15186 21437 15219 21439
rect 6814 21129 6847 21130
rect 11092 21129 11125 21130
rect 12380 21129 12413 21130
rect 12932 21129 12965 21130
rect 6814 21128 12965 21129
rect 6814 21100 6817 21128
rect 6845 21100 11095 21128
rect 11123 21100 12383 21128
rect 12411 21100 12935 21128
rect 12963 21100 12965 21128
rect 6814 21099 12965 21100
rect 6814 21097 6847 21099
rect 11092 21097 11125 21099
rect 12380 21097 12413 21099
rect 12932 21097 12965 21099
rect 11138 20857 11171 20858
rect 11276 20857 11309 20858
rect 11138 20856 11309 20857
rect 11138 20828 11141 20856
rect 11169 20828 11279 20856
rect 11307 20828 11309 20856
rect 11138 20827 11309 20828
rect 11138 20825 11171 20827
rect 11276 20825 11309 20827
rect 5756 20789 5789 20790
rect 5848 20789 5881 20790
rect 10218 20789 10251 20790
rect 5756 20788 10251 20789
rect 5756 20760 5759 20788
rect 5787 20760 5851 20788
rect 5879 20760 10221 20788
rect 10249 20760 10251 20788
rect 5756 20759 10251 20760
rect 5756 20757 5789 20759
rect 5848 20757 5881 20759
rect 10218 20757 10251 20759
rect 12380 20245 12413 20246
rect 14082 20245 14115 20246
rect 14404 20245 14437 20246
rect 12380 20244 14437 20245
rect 12380 20216 12383 20244
rect 12411 20216 14085 20244
rect 14113 20216 14407 20244
rect 14435 20216 14437 20244
rect 12380 20215 14437 20216
rect 12380 20213 12413 20215
rect 14082 20213 14115 20215
rect 14404 20213 14437 20215
rect 11920 20041 11953 20042
rect 14220 20041 14253 20042
rect 11920 20040 14253 20041
rect 11920 20012 11923 20040
rect 11951 20012 14223 20040
rect 14251 20012 14253 20040
rect 11920 20011 14253 20012
rect 11920 20009 11953 20011
rect 14220 20009 14253 20011
rect 12610 19973 12643 19974
rect 13116 19973 13149 19974
rect 12610 19972 13149 19973
rect 12610 19944 12613 19972
rect 12641 19944 13119 19972
rect 13147 19944 13149 19972
rect 12610 19943 13149 19944
rect 12610 19941 12643 19943
rect 13116 19941 13149 19943
rect 20752 19973 20785 19974
rect 22914 19973 22947 19974
rect 20752 19972 22947 19973
rect 20752 19944 20755 19972
rect 20783 19944 22917 19972
rect 22945 19944 22947 19972
rect 20752 19943 22947 19944
rect 20752 19941 20785 19943
rect 22914 19941 22947 19943
rect 6998 19701 7031 19702
rect 8700 19701 8733 19702
rect 11184 19701 11217 19702
rect 6998 19700 11217 19701
rect 6998 19672 7001 19700
rect 7029 19672 8703 19700
rect 8731 19672 11187 19700
rect 11215 19672 11217 19700
rect 6998 19671 11217 19672
rect 6998 19669 7031 19671
rect 8700 19669 8733 19671
rect 11184 19669 11217 19671
rect 22914 19565 22947 19566
rect 24386 19565 24419 19566
rect 22914 19564 24419 19565
rect 22914 19536 22917 19564
rect 22945 19536 24389 19564
rect 24417 19536 24419 19564
rect 22914 19535 24419 19536
rect 22914 19533 22947 19535
rect 24386 19533 24419 19535
rect 4928 19429 4961 19430
rect 5526 19429 5559 19430
rect 4928 19428 5559 19429
rect 4928 19400 4931 19428
rect 4959 19400 5529 19428
rect 5557 19400 5559 19428
rect 4928 19399 5559 19400
rect 4928 19397 4961 19399
rect 5526 19397 5559 19399
rect 10770 18613 10803 18614
rect 12656 18613 12689 18614
rect 10770 18612 12689 18613
rect 10770 18584 10773 18612
rect 10801 18584 12659 18612
rect 12687 18584 12689 18612
rect 10770 18583 12689 18584
rect 10770 18581 10803 18583
rect 12656 18581 12689 18583
rect 13116 18613 13149 18614
rect 14910 18613 14943 18614
rect 13116 18612 14943 18613
rect 13116 18584 13119 18612
rect 13147 18584 14913 18612
rect 14941 18584 14943 18612
rect 13116 18583 14943 18584
rect 13116 18581 13149 18583
rect 14910 18581 14943 18583
rect 21626 18613 21659 18614
rect 24478 18613 24511 18614
rect 21626 18612 24511 18613
rect 21626 18584 21629 18612
rect 21657 18584 24481 18612
rect 24509 18584 24511 18612
rect 21626 18583 24511 18584
rect 21626 18581 21659 18583
rect 24478 18581 24511 18583
rect 4836 18545 4869 18546
rect 0 18544 4869 18545
rect 0 18516 4839 18544
rect 4867 18516 4869 18544
rect 0 18515 4869 18516
rect 4836 18513 4869 18515
rect 20338 18545 20371 18546
rect 20614 18545 20647 18546
rect 22454 18545 22487 18546
rect 20338 18544 22487 18545
rect 20338 18516 20341 18544
rect 20369 18516 20617 18544
rect 20645 18516 22457 18544
rect 22485 18516 22487 18544
rect 20338 18515 22487 18516
rect 20338 18513 20371 18515
rect 20614 18513 20647 18515
rect 22454 18513 22487 18515
rect 18682 18477 18715 18478
rect 18912 18477 18945 18478
rect 23052 18477 23085 18478
rect 18682 18476 23085 18477
rect 18682 18448 18685 18476
rect 18713 18448 18915 18476
rect 18943 18448 23055 18476
rect 23083 18448 23085 18476
rect 18682 18447 23085 18448
rect 18682 18445 18715 18447
rect 18912 18445 18945 18447
rect 23052 18445 23085 18447
rect 5020 18409 5053 18410
rect 9528 18409 9561 18410
rect 10816 18409 10849 18410
rect 5020 18408 10849 18409
rect 5020 18380 5023 18408
rect 5051 18380 9531 18408
rect 9559 18380 10819 18408
rect 10847 18380 10849 18408
rect 5020 18379 10849 18380
rect 5020 18377 5053 18379
rect 9528 18377 9561 18379
rect 10816 18377 10849 18379
rect 20936 18409 20969 18410
rect 24478 18409 24511 18410
rect 20936 18408 24511 18409
rect 20936 18380 20939 18408
rect 20967 18380 24481 18408
rect 24509 18380 24511 18408
rect 20936 18379 24511 18380
rect 20936 18377 20969 18379
rect 24478 18377 24511 18379
rect 13622 18137 13655 18138
rect 14588 18137 14621 18138
rect 13622 18136 14621 18137
rect 13622 18108 13625 18136
rect 13653 18108 14591 18136
rect 14619 18108 14621 18136
rect 13622 18107 14621 18108
rect 13622 18105 13655 18107
rect 14588 18105 14621 18107
rect 22040 17525 22073 17526
rect 23972 17525 24005 17526
rect 22040 17524 24005 17525
rect 22040 17496 22043 17524
rect 22071 17496 23975 17524
rect 24003 17496 24005 17524
rect 22040 17495 24005 17496
rect 22040 17493 22073 17495
rect 23972 17493 24005 17495
rect 23236 17389 23269 17390
rect 25582 17389 25615 17390
rect 25904 17389 25937 17390
rect 23236 17388 25937 17389
rect 23236 17360 23239 17388
rect 23267 17360 25585 17388
rect 25613 17360 25907 17388
rect 25935 17360 25937 17388
rect 23236 17359 25937 17360
rect 23236 17357 23269 17359
rect 25582 17357 25615 17359
rect 25904 17357 25937 17359
rect 12886 17049 12919 17050
rect 12886 17048 15885 17049
rect 12886 17020 12889 17048
rect 12917 17020 15885 17048
rect 12886 17019 15885 17020
rect 12886 17017 12919 17019
rect 12242 16981 12275 16982
rect 15140 16981 15173 16982
rect 12242 16980 15173 16981
rect 12242 16952 12245 16980
rect 12273 16952 15143 16980
rect 15171 16952 15173 16980
rect 12242 16951 15173 16952
rect 15855 16981 15885 17019
rect 16014 16981 16047 16982
rect 16474 16981 16507 16982
rect 15855 16980 16507 16981
rect 15855 16952 16017 16980
rect 16045 16952 16477 16980
rect 16505 16952 16507 16980
rect 15855 16951 16507 16952
rect 12242 16949 12275 16951
rect 15140 16949 15173 16951
rect 16014 16949 16047 16951
rect 16474 16949 16507 16951
rect 20108 16913 20141 16914
rect 22684 16913 22717 16914
rect 20108 16912 22717 16913
rect 20108 16884 20111 16912
rect 20139 16884 22687 16912
rect 22715 16884 22717 16912
rect 20108 16883 22717 16884
rect 20108 16881 20141 16883
rect 22684 16881 22717 16883
rect 13162 16845 13195 16846
rect 15554 16845 15587 16846
rect 13162 16844 15587 16845
rect 13162 16816 13165 16844
rect 13193 16816 15557 16844
rect 15585 16816 15587 16844
rect 13162 16815 15587 16816
rect 13162 16813 13195 16815
rect 15554 16813 15587 16815
rect 11736 16777 11769 16778
rect 14634 16777 14667 16778
rect 11736 16776 14667 16777
rect 11736 16748 11739 16776
rect 11767 16748 14637 16776
rect 14665 16748 14667 16776
rect 11736 16747 14667 16748
rect 11736 16745 11769 16747
rect 14634 16745 14667 16747
rect 15508 16777 15541 16778
rect 15968 16777 16001 16778
rect 15508 16776 16001 16777
rect 15508 16748 15511 16776
rect 15539 16748 15971 16776
rect 15999 16748 16001 16776
rect 15508 16747 16001 16748
rect 15508 16745 15541 16747
rect 15968 16745 16001 16747
rect 14542 16709 14575 16710
rect 17118 16709 17151 16710
rect 14542 16708 17151 16709
rect 14542 16680 14545 16708
rect 14573 16680 17121 16708
rect 17149 16680 17151 16708
rect 14542 16679 17151 16680
rect 14542 16677 14575 16679
rect 17118 16677 17151 16679
rect 21258 16641 21291 16642
rect 21350 16641 21383 16642
rect 26134 16641 26167 16642
rect 21258 16640 26167 16641
rect 21258 16612 21261 16640
rect 21289 16612 21353 16640
rect 21381 16612 26137 16640
rect 26165 16612 26167 16640
rect 21258 16611 26167 16612
rect 21258 16609 21291 16611
rect 21350 16609 21383 16611
rect 26134 16609 26167 16611
rect 4744 16437 4777 16438
rect 6768 16437 6801 16438
rect 4744 16436 6801 16437
rect 4744 16408 4747 16436
rect 4775 16408 6771 16436
rect 6799 16408 6801 16436
rect 4744 16407 6801 16408
rect 4744 16405 4777 16407
rect 6768 16405 6801 16407
rect 4284 16301 4317 16302
rect 4928 16301 4961 16302
rect 4284 16300 4961 16301
rect 4284 16272 4287 16300
rect 4315 16272 4931 16300
rect 4959 16272 4961 16300
rect 4284 16271 4961 16272
rect 4284 16269 4317 16271
rect 4928 16269 4961 16271
rect 5986 16301 6019 16302
rect 9022 16301 9055 16302
rect 11184 16301 11217 16302
rect 5986 16300 11217 16301
rect 5986 16272 5989 16300
rect 6017 16272 9025 16300
rect 9053 16272 11187 16300
rect 11215 16272 11217 16300
rect 5986 16271 11217 16272
rect 5986 16269 6019 16271
rect 9022 16269 9055 16271
rect 11184 16269 11217 16271
rect 3134 16233 3167 16234
rect 4514 16233 4547 16234
rect 3134 16232 4547 16233
rect 3134 16204 3137 16232
rect 3165 16204 4517 16232
rect 4545 16204 4547 16232
rect 3134 16203 4547 16204
rect 3134 16201 3167 16203
rect 4514 16201 4547 16203
rect 18636 15757 18669 15758
rect 20982 15757 21015 15758
rect 18636 15756 21015 15757
rect 18636 15728 18639 15756
rect 18667 15728 20985 15756
rect 21013 15728 21015 15756
rect 18636 15727 21015 15728
rect 18636 15725 18669 15727
rect 20982 15725 21015 15727
rect 27560 15281 27593 15282
rect 29722 15281 29755 15282
rect 27560 15280 29755 15281
rect 27560 15252 27563 15280
rect 27591 15252 29725 15280
rect 29753 15252 29755 15280
rect 27560 15251 29755 15252
rect 27560 15249 27593 15251
rect 29722 15249 29755 15251
rect 31746 15281 31779 15282
rect 31746 15280 33000 15281
rect 31746 15252 31749 15280
rect 31777 15252 33000 15280
rect 31746 15251 33000 15252
rect 31746 15249 31779 15251
rect 26962 15213 26995 15214
rect 28342 15213 28375 15214
rect 26962 15212 28375 15213
rect 26962 15184 26965 15212
rect 26993 15184 28345 15212
rect 28373 15184 28375 15212
rect 26962 15183 28375 15184
rect 26962 15181 26995 15183
rect 28342 15181 28375 15183
rect 7136 15145 7169 15146
rect 7596 15145 7629 15146
rect 7136 15144 7629 15145
rect 7136 15116 7139 15144
rect 7167 15116 7599 15144
rect 7627 15116 7629 15144
rect 7136 15115 7629 15116
rect 7136 15113 7169 15115
rect 7596 15113 7629 15115
rect 12104 15145 12137 15146
rect 14542 15145 14575 15146
rect 12104 15144 14575 15145
rect 12104 15116 12107 15144
rect 12135 15116 14545 15144
rect 14573 15116 14575 15144
rect 12104 15115 14575 15116
rect 12104 15113 12137 15115
rect 14542 15113 14575 15115
rect 6032 14601 6065 14602
rect 6814 14601 6847 14602
rect 7780 14601 7813 14602
rect 6032 14600 7813 14601
rect 6032 14572 6035 14600
rect 6063 14572 6817 14600
rect 6845 14572 7783 14600
rect 7811 14572 7813 14600
rect 6032 14571 7813 14572
rect 6032 14569 6065 14571
rect 6814 14569 6847 14571
rect 7780 14569 7813 14571
rect 4882 14533 4915 14534
rect 7918 14533 7951 14534
rect 4882 14532 7951 14533
rect 4882 14504 4885 14532
rect 4913 14504 7921 14532
rect 7949 14504 7951 14532
rect 4882 14503 7951 14504
rect 4882 14501 4915 14503
rect 7918 14501 7951 14503
rect 12380 14533 12413 14534
rect 13254 14533 13287 14534
rect 12380 14532 13287 14533
rect 12380 14504 12383 14532
rect 12411 14504 13257 14532
rect 13285 14504 13287 14532
rect 12380 14503 13287 14504
rect 12380 14501 12413 14503
rect 13254 14501 13287 14503
rect 8746 13717 8779 13718
rect 10908 13717 10941 13718
rect 14036 13717 14069 13718
rect 14542 13717 14575 13718
rect 8746 13716 14575 13717
rect 8746 13688 8749 13716
rect 8777 13688 10911 13716
rect 10939 13688 14039 13716
rect 14067 13688 14545 13716
rect 14573 13688 14575 13716
rect 8746 13687 14575 13688
rect 8746 13685 8779 13687
rect 10908 13685 10941 13687
rect 14036 13685 14069 13687
rect 14542 13685 14575 13687
rect 14128 13649 14161 13650
rect 16290 13649 16323 13650
rect 14128 13648 16323 13649
rect 14128 13620 14131 13648
rect 14159 13620 16293 13648
rect 16321 13620 16323 13648
rect 14128 13619 16323 13620
rect 14128 13617 14161 13619
rect 16290 13617 16323 13619
rect 10264 13581 10297 13582
rect 14726 13581 14759 13582
rect 15370 13581 15403 13582
rect 10264 13580 15403 13581
rect 10264 13552 10267 13580
rect 10295 13552 14729 13580
rect 14757 13552 15373 13580
rect 15401 13552 15403 13580
rect 10264 13551 15403 13552
rect 10264 13549 10297 13551
rect 14726 13549 14759 13551
rect 15370 13549 15403 13551
rect 18314 13513 18347 13514
rect 19050 13513 19083 13514
rect 18314 13512 19083 13513
rect 18314 13484 18317 13512
rect 18345 13484 19053 13512
rect 19081 13484 19083 13512
rect 18314 13483 19083 13484
rect 18314 13481 18347 13483
rect 19050 13481 19083 13483
rect 8976 13377 9009 13378
rect 6195 13376 9009 13377
rect 6195 13348 8979 13376
rect 9007 13348 9009 13376
rect 6195 13347 9009 13348
rect 4744 13309 4777 13310
rect 6195 13309 6225 13347
rect 8976 13345 9009 13347
rect 4744 13308 6225 13309
rect 4744 13280 4747 13308
rect 4775 13280 6225 13308
rect 4744 13279 6225 13280
rect 7182 13309 7215 13310
rect 10080 13309 10113 13310
rect 7182 13308 10113 13309
rect 7182 13280 7185 13308
rect 7213 13280 10083 13308
rect 10111 13280 10113 13308
rect 7182 13279 10113 13280
rect 4744 13277 4777 13279
rect 7182 13277 7215 13279
rect 10080 13277 10113 13279
rect 11736 13309 11769 13310
rect 14956 13309 14989 13310
rect 11736 13308 14989 13309
rect 11736 13280 11739 13308
rect 11767 13280 14959 13308
rect 14987 13280 14989 13308
rect 11736 13279 14989 13280
rect 11736 13277 11769 13279
rect 14956 13277 14989 13279
rect 8194 13241 8227 13242
rect 12058 13241 12091 13242
rect 8194 13240 14505 13241
rect 8194 13212 8197 13240
rect 8225 13212 12061 13240
rect 12089 13212 14505 13240
rect 8194 13211 14505 13212
rect 8194 13209 8227 13211
rect 12058 13209 12091 13211
rect 8102 13173 8135 13174
rect 11736 13173 11769 13174
rect 8102 13172 11769 13173
rect 8102 13144 8105 13172
rect 8133 13144 11739 13172
rect 11767 13144 11769 13172
rect 8102 13143 11769 13144
rect 14475 13173 14505 13211
rect 14634 13173 14667 13174
rect 14475 13172 14667 13173
rect 14475 13144 14637 13172
rect 14665 13144 14667 13172
rect 14475 13143 14667 13144
rect 8102 13141 8135 13143
rect 11736 13141 11769 13143
rect 14634 13141 14667 13143
rect 19234 12969 19267 12970
rect 23926 12969 23959 12970
rect 19234 12968 23959 12969
rect 19234 12940 19237 12968
rect 19265 12940 23929 12968
rect 23957 12940 23959 12968
rect 19234 12939 23959 12940
rect 19234 12937 19267 12939
rect 23926 12937 23959 12939
rect 21626 12697 21659 12698
rect 24800 12697 24833 12698
rect 21626 12696 24833 12697
rect 21626 12668 21629 12696
rect 21657 12668 24803 12696
rect 24831 12668 24833 12696
rect 21626 12667 24833 12668
rect 21626 12665 21659 12667
rect 24800 12665 24833 12667
rect 3410 12629 3443 12630
rect 9022 12629 9055 12630
rect 3410 12628 9055 12629
rect 3410 12600 3413 12628
rect 3441 12600 9025 12628
rect 9053 12600 9055 12628
rect 3410 12599 9055 12600
rect 3410 12597 3443 12599
rect 9022 12597 9055 12599
rect 20430 12629 20463 12630
rect 26226 12629 26259 12630
rect 20430 12628 26259 12629
rect 20430 12600 20433 12628
rect 20461 12600 26229 12628
rect 26257 12600 26259 12628
rect 20430 12599 26259 12600
rect 20430 12597 20463 12599
rect 26226 12597 26259 12599
rect 6906 12493 6939 12494
rect 10402 12493 10435 12494
rect 6906 12492 10435 12493
rect 6906 12464 6909 12492
rect 6937 12464 10405 12492
rect 10433 12464 10435 12492
rect 6906 12463 10435 12464
rect 6906 12461 6939 12463
rect 10402 12461 10435 12463
rect 7596 12425 7629 12426
rect 7918 12425 7951 12426
rect 11644 12425 11677 12426
rect 13852 12425 13885 12426
rect 7596 12424 13885 12425
rect 7596 12396 7599 12424
rect 7627 12396 7921 12424
rect 7949 12396 11647 12424
rect 11675 12396 13855 12424
rect 13883 12396 13885 12424
rect 7596 12395 13885 12396
rect 7596 12393 7629 12395
rect 7918 12393 7951 12395
rect 11644 12393 11677 12395
rect 13852 12393 13885 12395
rect 13162 12357 13195 12358
rect 15278 12357 15311 12358
rect 13162 12356 15311 12357
rect 13162 12328 13165 12356
rect 13193 12328 15281 12356
rect 15309 12328 15311 12356
rect 13162 12327 15311 12328
rect 13162 12325 13195 12327
rect 15278 12325 15311 12327
rect 9666 12153 9699 12154
rect 12012 12153 12045 12154
rect 14496 12153 14529 12154
rect 9666 12152 14529 12153
rect 9666 12124 9669 12152
rect 9697 12124 12015 12152
rect 12043 12124 14499 12152
rect 14527 12124 14529 12152
rect 9666 12123 14529 12124
rect 9666 12121 9699 12123
rect 12012 12121 12045 12123
rect 14496 12121 14529 12123
rect 5388 12017 5421 12018
rect 0 12016 5421 12017
rect 0 11988 5391 12016
rect 5419 11988 5421 12016
rect 0 11987 5421 11988
rect 5388 11985 5421 11987
rect 7320 11949 7353 11950
rect 9988 11949 10021 11950
rect 7320 11948 10021 11949
rect 7320 11920 7323 11948
rect 7351 11920 9991 11948
rect 10019 11920 10021 11948
rect 7320 11919 10021 11920
rect 7320 11917 7353 11919
rect 9988 11917 10021 11919
rect 13024 11949 13057 11950
rect 15462 11949 15495 11950
rect 13024 11948 15495 11949
rect 13024 11920 13027 11948
rect 13055 11920 15465 11948
rect 15493 11920 15495 11948
rect 13024 11919 15495 11920
rect 13024 11917 13057 11919
rect 15462 11917 15495 11919
rect 9114 11881 9147 11882
rect 11736 11881 11769 11882
rect 14404 11881 14437 11882
rect 9114 11880 14437 11881
rect 9114 11852 9117 11880
rect 9145 11852 11739 11880
rect 11767 11852 14407 11880
rect 14435 11852 14437 11880
rect 9114 11851 14437 11852
rect 9114 11849 9147 11851
rect 11736 11849 11769 11851
rect 14404 11849 14437 11851
rect 8792 11813 8825 11814
rect 11046 11813 11079 11814
rect 11644 11813 11677 11814
rect 8792 11812 11677 11813
rect 8792 11784 8795 11812
rect 8823 11784 11049 11812
rect 11077 11784 11647 11812
rect 11675 11784 11677 11812
rect 8792 11783 11677 11784
rect 8792 11781 8825 11783
rect 11046 11781 11079 11783
rect 11644 11781 11677 11783
rect 9574 11745 9607 11746
rect 11920 11745 11953 11746
rect 14358 11745 14391 11746
rect 9574 11744 14391 11745
rect 9574 11716 9577 11744
rect 9605 11716 11923 11744
rect 11951 11716 14361 11744
rect 14389 11716 14391 11744
rect 9574 11715 14391 11716
rect 9574 11713 9607 11715
rect 11920 11713 11953 11715
rect 14358 11713 14391 11715
rect 26180 11745 26213 11746
rect 28204 11745 28237 11746
rect 26180 11744 28237 11745
rect 26180 11716 26183 11744
rect 26211 11716 28207 11744
rect 28235 11716 28237 11744
rect 26180 11715 28237 11716
rect 26180 11713 26213 11715
rect 28204 11713 28237 11715
rect 6860 11473 6893 11474
rect 8700 11473 8733 11474
rect 6860 11472 8733 11473
rect 6860 11444 6863 11472
rect 6891 11444 8703 11472
rect 8731 11444 8733 11472
rect 6860 11443 8733 11444
rect 6860 11441 6893 11443
rect 8700 11441 8733 11443
rect 21350 10861 21383 10862
rect 23512 10861 23545 10862
rect 21350 10860 23545 10861
rect 21350 10832 21353 10860
rect 21381 10832 23515 10860
rect 23543 10832 23545 10860
rect 21350 10831 23545 10832
rect 21350 10829 21383 10831
rect 23512 10829 23545 10831
rect 22914 10793 22947 10794
rect 23374 10793 23407 10794
rect 22914 10792 33000 10793
rect 22914 10764 22917 10792
rect 22945 10764 23377 10792
rect 23405 10764 33000 10792
rect 22914 10763 33000 10764
rect 22914 10761 22947 10763
rect 23374 10761 23407 10763
rect 25582 10725 25615 10726
rect 27744 10725 27777 10726
rect 25582 10724 27777 10725
rect 25582 10696 25585 10724
rect 25613 10696 27747 10724
rect 27775 10696 27777 10724
rect 25582 10695 27777 10696
rect 25582 10693 25615 10695
rect 27744 10693 27777 10695
rect 22684 10453 22717 10454
rect 23420 10453 23453 10454
rect 26226 10453 26259 10454
rect 22684 10452 26259 10453
rect 22684 10424 22687 10452
rect 22715 10424 23423 10452
rect 23451 10424 26229 10452
rect 26257 10424 26259 10452
rect 22684 10423 26259 10424
rect 22684 10421 22717 10423
rect 23420 10421 23453 10423
rect 26226 10421 26259 10423
rect 16771 10354 16774 10386
rect 16806 10385 16809 10386
rect 17072 10385 17105 10386
rect 16806 10384 17105 10385
rect 16806 10356 17075 10384
rect 17103 10356 17105 10384
rect 16806 10355 17105 10356
rect 16806 10354 16809 10355
rect 17072 10353 17105 10355
rect 16704 9637 16737 9638
rect 16771 9637 16774 9638
rect 16704 9636 16774 9637
rect 16704 9608 16707 9636
rect 16735 9608 16774 9636
rect 16704 9607 16774 9608
rect 16704 9605 16737 9607
rect 16771 9606 16774 9607
rect 16806 9606 16809 9638
rect 20430 9501 20463 9502
rect 28802 9501 28835 9502
rect 29676 9501 29709 9502
rect 20430 9500 29709 9501
rect 20430 9472 20433 9500
rect 20461 9472 28805 9500
rect 28833 9472 29679 9500
rect 29707 9472 29709 9500
rect 20430 9471 29709 9472
rect 20430 9469 20463 9471
rect 28802 9469 28835 9471
rect 29676 9469 29709 9471
rect 26686 9433 26719 9434
rect 28020 9433 28053 9434
rect 28388 9433 28421 9434
rect 26686 9432 28421 9433
rect 26686 9404 26689 9432
rect 26717 9404 28023 9432
rect 28051 9404 28391 9432
rect 28419 9404 28421 9432
rect 26686 9403 28421 9404
rect 26686 9401 26719 9403
rect 28020 9401 28053 9403
rect 28388 9401 28421 9403
rect 22408 9365 22441 9366
rect 22960 9365 22993 9366
rect 26962 9365 26995 9366
rect 22408 9364 26995 9365
rect 22408 9336 22411 9364
rect 22439 9336 22963 9364
rect 22991 9336 26965 9364
rect 26993 9336 26995 9364
rect 22408 9335 26995 9336
rect 22408 9333 22441 9335
rect 22960 9333 22993 9335
rect 26962 9333 26995 9335
rect 21350 9297 21383 9298
rect 25352 9297 25385 9298
rect 21350 9296 25385 9297
rect 21350 9268 21353 9296
rect 21381 9268 25355 9296
rect 25383 9268 25385 9296
rect 21350 9267 25385 9268
rect 21350 9265 21383 9267
rect 25352 9265 25385 9267
rect 20936 9229 20969 9230
rect 25858 9229 25891 9230
rect 20936 9228 25891 9229
rect 20936 9200 20939 9228
rect 20967 9200 25861 9228
rect 25889 9200 25891 9228
rect 20936 9199 25891 9200
rect 20936 9197 20969 9199
rect 25858 9197 25891 9199
rect 28066 9229 28099 9230
rect 28296 9229 28329 9230
rect 28066 9228 28329 9229
rect 28066 9200 28069 9228
rect 28097 9200 28299 9228
rect 28327 9200 28329 9228
rect 28066 9199 28329 9200
rect 28066 9197 28099 9199
rect 28296 9197 28329 9199
rect 23880 9161 23913 9162
rect 25720 9161 25753 9162
rect 23880 9160 25753 9161
rect 23880 9132 23883 9160
rect 23911 9132 25723 9160
rect 25751 9132 25753 9160
rect 23880 9131 25753 9132
rect 23880 9129 23913 9131
rect 25720 9129 25753 9131
rect 24202 9025 24235 9026
rect 28066 9025 28099 9026
rect 24202 9024 28099 9025
rect 24202 8996 24205 9024
rect 24233 8996 28069 9024
rect 28097 8996 28099 9024
rect 24202 8995 28099 8996
rect 24202 8993 24235 8995
rect 28066 8993 28099 8995
rect 24616 8277 24649 8278
rect 29722 8277 29755 8278
rect 24616 8276 29755 8277
rect 24616 8248 24619 8276
rect 24647 8248 29725 8276
rect 29753 8248 29755 8276
rect 24616 8247 29755 8248
rect 24616 8245 24649 8247
rect 29722 8245 29755 8247
rect 8746 7665 8770 7666
rect 8724 7664 8770 7665
rect 8724 7636 8749 7664
rect 8724 7635 8770 7636
rect 8746 7634 8770 7635
rect 8802 7634 8805 7666
rect 8746 7633 8779 7634
rect 7136 7597 7169 7598
rect 8838 7597 8871 7598
rect 7136 7596 8871 7597
rect 7136 7568 7139 7596
rect 7167 7568 8841 7596
rect 8869 7568 8871 7596
rect 7136 7567 8871 7568
rect 7136 7565 7169 7567
rect 8838 7565 8871 7567
rect 23512 7597 23545 7598
rect 28572 7597 28605 7598
rect 23512 7596 28605 7597
rect 23512 7568 23515 7596
rect 23543 7568 28575 7596
rect 28603 7568 28605 7596
rect 23512 7567 28605 7568
rect 23512 7565 23545 7567
rect 28572 7565 28605 7567
rect 24202 7189 24235 7190
rect 27882 7189 27915 7190
rect 24202 7188 27915 7189
rect 24202 7160 24205 7188
rect 24233 7160 27885 7188
rect 27913 7160 27915 7188
rect 24202 7159 27915 7160
rect 24202 7157 24235 7159
rect 27882 7157 27915 7159
rect 24892 7053 24925 7054
rect 28894 7053 28927 7054
rect 24892 7052 28927 7053
rect 24892 7024 24895 7052
rect 24923 7024 28897 7052
rect 28925 7024 28927 7052
rect 24892 7023 28927 7024
rect 24892 7021 24925 7023
rect 28894 7021 28927 7023
rect 21948 6985 21981 6986
rect 29124 6985 29157 6986
rect 21948 6984 29157 6985
rect 21948 6956 21951 6984
rect 21979 6956 29127 6984
rect 29155 6956 29157 6984
rect 21948 6955 29157 6956
rect 21948 6953 21981 6955
rect 29124 6953 29157 6955
rect 22592 6917 22625 6918
rect 27100 6917 27133 6918
rect 22592 6916 27133 6917
rect 22592 6888 22595 6916
rect 22623 6888 27103 6916
rect 27131 6888 27133 6916
rect 22592 6887 27133 6888
rect 22592 6885 22625 6887
rect 27100 6885 27133 6887
rect 20568 6849 20601 6850
rect 23512 6849 23545 6850
rect 20568 6848 23545 6849
rect 20568 6820 20571 6848
rect 20599 6820 23515 6848
rect 23543 6820 23545 6848
rect 20568 6819 23545 6820
rect 20568 6817 20601 6819
rect 23512 6817 23545 6819
rect 21258 6713 21291 6714
rect 28204 6713 28237 6714
rect 21258 6712 28237 6713
rect 21258 6684 21261 6712
rect 21289 6684 28207 6712
rect 28235 6684 28237 6712
rect 21258 6683 28237 6684
rect 21258 6681 21291 6683
rect 28204 6681 28237 6683
rect 26226 6645 26259 6646
rect 26962 6645 26995 6646
rect 26159 6644 26995 6645
rect 26159 6616 26229 6644
rect 26257 6616 26965 6644
rect 26993 6616 26995 6644
rect 26159 6615 26995 6616
rect 21442 6577 21475 6578
rect 26159 6577 26189 6615
rect 26226 6613 26259 6615
rect 26962 6613 26995 6615
rect 21442 6576 26189 6577
rect 21442 6548 21445 6576
rect 21473 6548 26189 6576
rect 21442 6547 26189 6548
rect 21442 6545 21475 6547
rect 21304 6509 21337 6510
rect 23420 6509 23453 6510
rect 28480 6509 28513 6510
rect 21304 6508 28513 6509
rect 21304 6480 21307 6508
rect 21335 6480 23423 6508
rect 23451 6480 28483 6508
rect 28511 6480 28513 6508
rect 21304 6479 28513 6480
rect 21304 6477 21337 6479
rect 23420 6477 23453 6479
rect 28480 6477 28513 6479
rect 5204 5625 5237 5626
rect 0 5624 5237 5625
rect 0 5596 5207 5624
rect 5235 5596 5237 5624
rect 0 5595 5237 5596
rect 5204 5593 5237 5595
rect 21442 5013 21475 5014
rect 24202 5013 24235 5014
rect 25858 5013 25891 5014
rect 21442 5012 25891 5013
rect 21442 4984 21445 5012
rect 21473 4984 24205 5012
rect 24233 4984 25861 5012
rect 25889 4984 25891 5012
rect 21442 4983 25891 4984
rect 21442 4981 21475 4983
rect 24202 4981 24235 4983
rect 25858 4981 25891 4983
rect 5526 661 5559 662
rect 8767 661 8770 662
rect 5526 660 8770 661
rect 5526 632 5529 660
rect 5557 632 8770 660
rect 5526 631 8770 632
rect 5526 629 5559 631
rect 8767 630 8770 631
rect 8802 630 8805 662
<< via3 >>
rect 16774 10354 16806 10386
rect 16774 9606 16806 9638
rect 8770 7664 8802 7666
rect 8770 7636 8777 7664
rect 8777 7636 8802 7664
rect 8770 7634 8802 7636
rect 8770 630 8802 662
<< metal4 >>
rect 4956 29323 5116 29344
rect 4956 29205 4977 29323
rect 5095 29205 5116 29323
rect 3956 28323 4116 28344
rect 3956 28205 3977 28323
rect 4095 28205 4116 28323
rect 3956 26323 4116 28205
rect 3956 26205 3977 26323
rect 4095 26205 4116 26323
rect 3956 24323 4116 26205
rect 3956 24205 3977 24323
rect 4095 24205 4116 24323
rect 3956 22323 4116 24205
rect 3956 22205 3977 22323
rect 4095 22205 4116 22323
rect 3956 20323 4116 22205
rect 3956 20205 3977 20323
rect 4095 20205 4116 20323
rect 3956 18323 4116 20205
rect 3956 18205 3977 18323
rect 4095 18205 4116 18323
rect 3956 16323 4116 18205
rect 3956 16205 3977 16323
rect 4095 16205 4116 16323
rect 3956 14323 4116 16205
rect 3956 14205 3977 14323
rect 4095 14205 4116 14323
rect 3956 12323 4116 14205
rect 3956 12205 3977 12323
rect 4095 12205 4116 12323
rect 3956 10323 4116 12205
rect 3956 10205 3977 10323
rect 4095 10205 4116 10323
rect 3956 8323 4116 10205
rect 3956 8205 3977 8323
rect 4095 8205 4116 8323
rect 3956 6323 4116 8205
rect 3956 6205 3977 6323
rect 4095 6205 4116 6323
rect 3956 4323 4116 6205
rect 4956 27323 5116 29205
rect 6956 29323 7116 29344
rect 6956 29205 6977 29323
rect 7095 29205 7116 29323
rect 4956 27205 4977 27323
rect 5095 27205 5116 27323
rect 4956 25323 5116 27205
rect 4956 25205 4977 25323
rect 5095 25205 5116 25323
rect 4956 23323 5116 25205
rect 4956 23205 4977 23323
rect 5095 23205 5116 23323
rect 4956 21323 5116 23205
rect 4956 21205 4977 21323
rect 5095 21205 5116 21323
rect 4956 19323 5116 21205
rect 4956 19205 4977 19323
rect 5095 19205 5116 19323
rect 4956 17323 5116 19205
rect 4956 17205 4977 17323
rect 5095 17205 5116 17323
rect 4956 15323 5116 17205
rect 4956 15205 4977 15323
rect 5095 15205 5116 15323
rect 4956 13323 5116 15205
rect 4956 13205 4977 13323
rect 5095 13205 5116 13323
rect 4956 11323 5116 13205
rect 4956 11205 4977 11323
rect 5095 11205 5116 11323
rect 4956 9323 5116 11205
rect 4956 9205 4977 9323
rect 5095 9205 5116 9323
rect 4956 7323 5116 9205
rect 4956 7205 4977 7323
rect 5095 7205 5116 7323
rect 4956 5323 5116 7205
rect 4956 5205 4977 5323
rect 5095 5205 5116 5323
rect 4956 5184 5116 5205
rect 5956 28323 6116 28344
rect 5956 28205 5977 28323
rect 6095 28205 6116 28323
rect 5956 26323 6116 28205
rect 5956 26205 5977 26323
rect 6095 26205 6116 26323
rect 5956 24323 6116 26205
rect 5956 24205 5977 24323
rect 6095 24205 6116 24323
rect 5956 22323 6116 24205
rect 5956 22205 5977 22323
rect 6095 22205 6116 22323
rect 5956 20323 6116 22205
rect 5956 20205 5977 20323
rect 6095 20205 6116 20323
rect 5956 18323 6116 20205
rect 5956 18205 5977 18323
rect 6095 18205 6116 18323
rect 5956 16323 6116 18205
rect 5956 16205 5977 16323
rect 6095 16205 6116 16323
rect 5956 14323 6116 16205
rect 5956 14205 5977 14323
rect 6095 14205 6116 14323
rect 5956 12323 6116 14205
rect 5956 12205 5977 12323
rect 6095 12205 6116 12323
rect 5956 10323 6116 12205
rect 5956 10205 5977 10323
rect 6095 10205 6116 10323
rect 5956 8323 6116 10205
rect 5956 8205 5977 8323
rect 6095 8205 6116 8323
rect 5956 6323 6116 8205
rect 5956 6205 5977 6323
rect 6095 6205 6116 6323
rect 3956 4205 3977 4323
rect 4095 4205 4116 4323
rect 3956 4184 4116 4205
rect 5956 4323 6116 6205
rect 6956 27323 7116 29205
rect 8956 29323 9116 29344
rect 8956 29205 8977 29323
rect 9095 29205 9116 29323
rect 6956 27205 6977 27323
rect 7095 27205 7116 27323
rect 6956 25323 7116 27205
rect 6956 25205 6977 25323
rect 7095 25205 7116 25323
rect 6956 23323 7116 25205
rect 6956 23205 6977 23323
rect 7095 23205 7116 23323
rect 6956 21323 7116 23205
rect 6956 21205 6977 21323
rect 7095 21205 7116 21323
rect 6956 19323 7116 21205
rect 6956 19205 6977 19323
rect 7095 19205 7116 19323
rect 6956 17323 7116 19205
rect 6956 17205 6977 17323
rect 7095 17205 7116 17323
rect 6956 15323 7116 17205
rect 6956 15205 6977 15323
rect 7095 15205 7116 15323
rect 6956 13323 7116 15205
rect 6956 13205 6977 13323
rect 7095 13205 7116 13323
rect 6956 11323 7116 13205
rect 6956 11205 6977 11323
rect 7095 11205 7116 11323
rect 6956 9323 7116 11205
rect 6956 9205 6977 9323
rect 7095 9205 7116 9323
rect 6956 7323 7116 9205
rect 6956 7205 6977 7323
rect 7095 7205 7116 7323
rect 6956 5323 7116 7205
rect 6956 5205 6977 5323
rect 7095 5205 7116 5323
rect 6956 5184 7116 5205
rect 7956 28323 8116 28344
rect 7956 28205 7977 28323
rect 8095 28205 8116 28323
rect 7956 26323 8116 28205
rect 7956 26205 7977 26323
rect 8095 26205 8116 26323
rect 7956 24323 8116 26205
rect 7956 24205 7977 24323
rect 8095 24205 8116 24323
rect 7956 22323 8116 24205
rect 7956 22205 7977 22323
rect 8095 22205 8116 22323
rect 7956 20323 8116 22205
rect 7956 20205 7977 20323
rect 8095 20205 8116 20323
rect 7956 18323 8116 20205
rect 7956 18205 7977 18323
rect 8095 18205 8116 18323
rect 7956 16323 8116 18205
rect 7956 16205 7977 16323
rect 8095 16205 8116 16323
rect 7956 14323 8116 16205
rect 7956 14205 7977 14323
rect 8095 14205 8116 14323
rect 7956 12323 8116 14205
rect 7956 12205 7977 12323
rect 8095 12205 8116 12323
rect 7956 10323 8116 12205
rect 7956 10205 7977 10323
rect 8095 10205 8116 10323
rect 7956 8323 8116 10205
rect 7956 8205 7977 8323
rect 8095 8205 8116 8323
rect 7956 6323 8116 8205
rect 8956 27323 9116 29205
rect 10956 29323 11116 29344
rect 10956 29205 10977 29323
rect 11095 29205 11116 29323
rect 8956 27205 8977 27323
rect 9095 27205 9116 27323
rect 8956 25323 9116 27205
rect 8956 25205 8977 25323
rect 9095 25205 9116 25323
rect 8956 23323 9116 25205
rect 8956 23205 8977 23323
rect 9095 23205 9116 23323
rect 8956 21323 9116 23205
rect 8956 21205 8977 21323
rect 9095 21205 9116 21323
rect 8956 19323 9116 21205
rect 8956 19205 8977 19323
rect 9095 19205 9116 19323
rect 8956 17323 9116 19205
rect 8956 17205 8977 17323
rect 9095 17205 9116 17323
rect 8956 15323 9116 17205
rect 8956 15205 8977 15323
rect 9095 15205 9116 15323
rect 8956 13323 9116 15205
rect 8956 13205 8977 13323
rect 9095 13205 9116 13323
rect 8956 11323 9116 13205
rect 8956 11205 8977 11323
rect 9095 11205 9116 11323
rect 8956 9323 9116 11205
rect 8956 9205 8977 9323
rect 9095 9205 9116 9323
rect 8769 7634 8770 7666
rect 8769 7633 8802 7634
rect 7956 6205 7977 6323
rect 8095 6205 8116 6323
rect 5956 4205 5977 4323
rect 6095 4205 6116 4323
rect 5956 4184 6116 4205
rect 7956 4323 8116 6205
rect 7956 4205 7977 4323
rect 8095 4205 8116 4323
rect 7956 4184 8116 4205
rect 8771 662 8801 7633
rect 8956 7323 9116 9205
rect 8956 7205 8977 7323
rect 9095 7205 9116 7323
rect 8956 5323 9116 7205
rect 8956 5205 8977 5323
rect 9095 5205 9116 5323
rect 8956 5184 9116 5205
rect 9956 28323 10116 28344
rect 9956 28205 9977 28323
rect 10095 28205 10116 28323
rect 9956 26323 10116 28205
rect 9956 26205 9977 26323
rect 10095 26205 10116 26323
rect 9956 24323 10116 26205
rect 9956 24205 9977 24323
rect 10095 24205 10116 24323
rect 9956 22323 10116 24205
rect 9956 22205 9977 22323
rect 10095 22205 10116 22323
rect 9956 20323 10116 22205
rect 9956 20205 9977 20323
rect 10095 20205 10116 20323
rect 9956 18323 10116 20205
rect 9956 18205 9977 18323
rect 10095 18205 10116 18323
rect 9956 16323 10116 18205
rect 9956 16205 9977 16323
rect 10095 16205 10116 16323
rect 9956 14323 10116 16205
rect 9956 14205 9977 14323
rect 10095 14205 10116 14323
rect 9956 12323 10116 14205
rect 9956 12205 9977 12323
rect 10095 12205 10116 12323
rect 9956 10323 10116 12205
rect 9956 10205 9977 10323
rect 10095 10205 10116 10323
rect 9956 8323 10116 10205
rect 9956 8205 9977 8323
rect 10095 8205 10116 8323
rect 9956 6323 10116 8205
rect 9956 6205 9977 6323
rect 10095 6205 10116 6323
rect 9956 4323 10116 6205
rect 10956 27323 11116 29205
rect 12956 29323 13116 29344
rect 12956 29205 12977 29323
rect 13095 29205 13116 29323
rect 10956 27205 10977 27323
rect 11095 27205 11116 27323
rect 10956 25323 11116 27205
rect 10956 25205 10977 25323
rect 11095 25205 11116 25323
rect 10956 23323 11116 25205
rect 10956 23205 10977 23323
rect 11095 23205 11116 23323
rect 10956 21323 11116 23205
rect 10956 21205 10977 21323
rect 11095 21205 11116 21323
rect 10956 19323 11116 21205
rect 10956 19205 10977 19323
rect 11095 19205 11116 19323
rect 10956 17323 11116 19205
rect 10956 17205 10977 17323
rect 11095 17205 11116 17323
rect 10956 15323 11116 17205
rect 10956 15205 10977 15323
rect 11095 15205 11116 15323
rect 10956 13323 11116 15205
rect 10956 13205 10977 13323
rect 11095 13205 11116 13323
rect 10956 11323 11116 13205
rect 10956 11205 10977 11323
rect 11095 11205 11116 11323
rect 10956 9323 11116 11205
rect 10956 9205 10977 9323
rect 11095 9205 11116 9323
rect 10956 7323 11116 9205
rect 10956 7205 10977 7323
rect 11095 7205 11116 7323
rect 10956 5323 11116 7205
rect 10956 5205 10977 5323
rect 11095 5205 11116 5323
rect 10956 5184 11116 5205
rect 11956 28323 12116 28344
rect 11956 28205 11977 28323
rect 12095 28205 12116 28323
rect 11956 26323 12116 28205
rect 11956 26205 11977 26323
rect 12095 26205 12116 26323
rect 11956 24323 12116 26205
rect 11956 24205 11977 24323
rect 12095 24205 12116 24323
rect 11956 22323 12116 24205
rect 11956 22205 11977 22323
rect 12095 22205 12116 22323
rect 11956 20323 12116 22205
rect 11956 20205 11977 20323
rect 12095 20205 12116 20323
rect 11956 18323 12116 20205
rect 11956 18205 11977 18323
rect 12095 18205 12116 18323
rect 11956 16323 12116 18205
rect 11956 16205 11977 16323
rect 12095 16205 12116 16323
rect 11956 14323 12116 16205
rect 11956 14205 11977 14323
rect 12095 14205 12116 14323
rect 11956 12323 12116 14205
rect 11956 12205 11977 12323
rect 12095 12205 12116 12323
rect 11956 10323 12116 12205
rect 11956 10205 11977 10323
rect 12095 10205 12116 10323
rect 11956 8323 12116 10205
rect 11956 8205 11977 8323
rect 12095 8205 12116 8323
rect 11956 6323 12116 8205
rect 11956 6205 11977 6323
rect 12095 6205 12116 6323
rect 9956 4205 9977 4323
rect 10095 4205 10116 4323
rect 9956 4184 10116 4205
rect 11956 4323 12116 6205
rect 12956 27323 13116 29205
rect 14956 29323 15116 29344
rect 14956 29205 14977 29323
rect 15095 29205 15116 29323
rect 12956 27205 12977 27323
rect 13095 27205 13116 27323
rect 12956 25323 13116 27205
rect 12956 25205 12977 25323
rect 13095 25205 13116 25323
rect 12956 23323 13116 25205
rect 12956 23205 12977 23323
rect 13095 23205 13116 23323
rect 12956 21323 13116 23205
rect 12956 21205 12977 21323
rect 13095 21205 13116 21323
rect 12956 19323 13116 21205
rect 12956 19205 12977 19323
rect 13095 19205 13116 19323
rect 12956 17323 13116 19205
rect 12956 17205 12977 17323
rect 13095 17205 13116 17323
rect 12956 15323 13116 17205
rect 12956 15205 12977 15323
rect 13095 15205 13116 15323
rect 12956 13323 13116 15205
rect 12956 13205 12977 13323
rect 13095 13205 13116 13323
rect 12956 11323 13116 13205
rect 12956 11205 12977 11323
rect 13095 11205 13116 11323
rect 12956 9323 13116 11205
rect 12956 9205 12977 9323
rect 13095 9205 13116 9323
rect 12956 7323 13116 9205
rect 12956 7205 12977 7323
rect 13095 7205 13116 7323
rect 12956 5323 13116 7205
rect 12956 5205 12977 5323
rect 13095 5205 13116 5323
rect 12956 5184 13116 5205
rect 13956 28323 14116 28344
rect 13956 28205 13977 28323
rect 14095 28205 14116 28323
rect 13956 26323 14116 28205
rect 13956 26205 13977 26323
rect 14095 26205 14116 26323
rect 13956 24323 14116 26205
rect 13956 24205 13977 24323
rect 14095 24205 14116 24323
rect 13956 22323 14116 24205
rect 13956 22205 13977 22323
rect 14095 22205 14116 22323
rect 13956 20323 14116 22205
rect 13956 20205 13977 20323
rect 14095 20205 14116 20323
rect 13956 18323 14116 20205
rect 13956 18205 13977 18323
rect 14095 18205 14116 18323
rect 13956 16323 14116 18205
rect 13956 16205 13977 16323
rect 14095 16205 14116 16323
rect 13956 14323 14116 16205
rect 13956 14205 13977 14323
rect 14095 14205 14116 14323
rect 13956 12323 14116 14205
rect 13956 12205 13977 12323
rect 14095 12205 14116 12323
rect 13956 10323 14116 12205
rect 13956 10205 13977 10323
rect 14095 10205 14116 10323
rect 13956 8323 14116 10205
rect 13956 8205 13977 8323
rect 14095 8205 14116 8323
rect 13956 6323 14116 8205
rect 13956 6205 13977 6323
rect 14095 6205 14116 6323
rect 11956 4205 11977 4323
rect 12095 4205 12116 4323
rect 11956 4184 12116 4205
rect 13956 4323 14116 6205
rect 14956 27323 15116 29205
rect 16956 29323 17116 29344
rect 16956 29205 16977 29323
rect 17095 29205 17116 29323
rect 14956 27205 14977 27323
rect 15095 27205 15116 27323
rect 14956 25323 15116 27205
rect 14956 25205 14977 25323
rect 15095 25205 15116 25323
rect 14956 23323 15116 25205
rect 14956 23205 14977 23323
rect 15095 23205 15116 23323
rect 14956 21323 15116 23205
rect 14956 21205 14977 21323
rect 15095 21205 15116 21323
rect 14956 19323 15116 21205
rect 14956 19205 14977 19323
rect 15095 19205 15116 19323
rect 14956 17323 15116 19205
rect 14956 17205 14977 17323
rect 15095 17205 15116 17323
rect 14956 15323 15116 17205
rect 14956 15205 14977 15323
rect 15095 15205 15116 15323
rect 14956 13323 15116 15205
rect 14956 13205 14977 13323
rect 15095 13205 15116 13323
rect 14956 11323 15116 13205
rect 14956 11205 14977 11323
rect 15095 11205 15116 11323
rect 14956 9323 15116 11205
rect 14956 9205 14977 9323
rect 15095 9205 15116 9323
rect 14956 7323 15116 9205
rect 14956 7205 14977 7323
rect 15095 7205 15116 7323
rect 14956 5323 15116 7205
rect 14956 5205 14977 5323
rect 15095 5205 15116 5323
rect 14956 5184 15116 5205
rect 15956 28323 16116 28344
rect 15956 28205 15977 28323
rect 16095 28205 16116 28323
rect 15956 26323 16116 28205
rect 15956 26205 15977 26323
rect 16095 26205 16116 26323
rect 15956 24323 16116 26205
rect 15956 24205 15977 24323
rect 16095 24205 16116 24323
rect 15956 22323 16116 24205
rect 15956 22205 15977 22323
rect 16095 22205 16116 22323
rect 15956 20323 16116 22205
rect 15956 20205 15977 20323
rect 16095 20205 16116 20323
rect 15956 18323 16116 20205
rect 15956 18205 15977 18323
rect 16095 18205 16116 18323
rect 15956 16323 16116 18205
rect 15956 16205 15977 16323
rect 16095 16205 16116 16323
rect 15956 14323 16116 16205
rect 15956 14205 15977 14323
rect 16095 14205 16116 14323
rect 15956 12323 16116 14205
rect 15956 12205 15977 12323
rect 16095 12205 16116 12323
rect 15956 10323 16116 12205
rect 16956 27323 17116 29205
rect 18956 29323 19116 29344
rect 18956 29205 18977 29323
rect 19095 29205 19116 29323
rect 16956 27205 16977 27323
rect 17095 27205 17116 27323
rect 16956 25323 17116 27205
rect 16956 25205 16977 25323
rect 17095 25205 17116 25323
rect 16956 23323 17116 25205
rect 16956 23205 16977 23323
rect 17095 23205 17116 23323
rect 16956 21323 17116 23205
rect 16956 21205 16977 21323
rect 17095 21205 17116 21323
rect 16956 19323 17116 21205
rect 16956 19205 16977 19323
rect 17095 19205 17116 19323
rect 16956 17323 17116 19205
rect 16956 17205 16977 17323
rect 17095 17205 17116 17323
rect 16956 15323 17116 17205
rect 16956 15205 16977 15323
rect 17095 15205 17116 15323
rect 16956 13323 17116 15205
rect 16956 13205 16977 13323
rect 17095 13205 17116 13323
rect 16956 11323 17116 13205
rect 16956 11205 16977 11323
rect 17095 11205 17116 11323
rect 16773 10354 16774 10386
rect 16773 10353 16806 10354
rect 15956 10205 15977 10323
rect 16095 10205 16116 10323
rect 15956 8323 16116 10205
rect 16775 9638 16805 10353
rect 16773 9606 16774 9638
rect 16773 9605 16806 9606
rect 15956 8205 15977 8323
rect 16095 8205 16116 8323
rect 15956 6323 16116 8205
rect 15956 6205 15977 6323
rect 16095 6205 16116 6323
rect 13956 4205 13977 4323
rect 14095 4205 14116 4323
rect 13956 4184 14116 4205
rect 15956 4323 16116 6205
rect 16956 9323 17116 11205
rect 16956 9205 16977 9323
rect 17095 9205 17116 9323
rect 16956 7323 17116 9205
rect 16956 7205 16977 7323
rect 17095 7205 17116 7323
rect 16956 5323 17116 7205
rect 16956 5205 16977 5323
rect 17095 5205 17116 5323
rect 16956 5184 17116 5205
rect 17956 28323 18116 28344
rect 17956 28205 17977 28323
rect 18095 28205 18116 28323
rect 17956 26323 18116 28205
rect 17956 26205 17977 26323
rect 18095 26205 18116 26323
rect 17956 24323 18116 26205
rect 17956 24205 17977 24323
rect 18095 24205 18116 24323
rect 17956 22323 18116 24205
rect 17956 22205 17977 22323
rect 18095 22205 18116 22323
rect 17956 20323 18116 22205
rect 17956 20205 17977 20323
rect 18095 20205 18116 20323
rect 17956 18323 18116 20205
rect 17956 18205 17977 18323
rect 18095 18205 18116 18323
rect 17956 16323 18116 18205
rect 17956 16205 17977 16323
rect 18095 16205 18116 16323
rect 17956 14323 18116 16205
rect 17956 14205 17977 14323
rect 18095 14205 18116 14323
rect 17956 12323 18116 14205
rect 17956 12205 17977 12323
rect 18095 12205 18116 12323
rect 17956 10323 18116 12205
rect 17956 10205 17977 10323
rect 18095 10205 18116 10323
rect 17956 8323 18116 10205
rect 17956 8205 17977 8323
rect 18095 8205 18116 8323
rect 17956 6323 18116 8205
rect 17956 6205 17977 6323
rect 18095 6205 18116 6323
rect 15956 4205 15977 4323
rect 16095 4205 16116 4323
rect 15956 4184 16116 4205
rect 17956 4323 18116 6205
rect 18956 27323 19116 29205
rect 20956 29323 21116 29344
rect 20956 29205 20977 29323
rect 21095 29205 21116 29323
rect 18956 27205 18977 27323
rect 19095 27205 19116 27323
rect 18956 25323 19116 27205
rect 18956 25205 18977 25323
rect 19095 25205 19116 25323
rect 18956 23323 19116 25205
rect 18956 23205 18977 23323
rect 19095 23205 19116 23323
rect 18956 21323 19116 23205
rect 18956 21205 18977 21323
rect 19095 21205 19116 21323
rect 18956 19323 19116 21205
rect 18956 19205 18977 19323
rect 19095 19205 19116 19323
rect 18956 17323 19116 19205
rect 18956 17205 18977 17323
rect 19095 17205 19116 17323
rect 18956 15323 19116 17205
rect 18956 15205 18977 15323
rect 19095 15205 19116 15323
rect 18956 13323 19116 15205
rect 18956 13205 18977 13323
rect 19095 13205 19116 13323
rect 18956 11323 19116 13205
rect 18956 11205 18977 11323
rect 19095 11205 19116 11323
rect 18956 9323 19116 11205
rect 18956 9205 18977 9323
rect 19095 9205 19116 9323
rect 18956 7323 19116 9205
rect 18956 7205 18977 7323
rect 19095 7205 19116 7323
rect 18956 5323 19116 7205
rect 18956 5205 18977 5323
rect 19095 5205 19116 5323
rect 18956 5184 19116 5205
rect 19956 28323 20116 28344
rect 19956 28205 19977 28323
rect 20095 28205 20116 28323
rect 19956 26323 20116 28205
rect 19956 26205 19977 26323
rect 20095 26205 20116 26323
rect 19956 24323 20116 26205
rect 19956 24205 19977 24323
rect 20095 24205 20116 24323
rect 19956 22323 20116 24205
rect 19956 22205 19977 22323
rect 20095 22205 20116 22323
rect 19956 20323 20116 22205
rect 19956 20205 19977 20323
rect 20095 20205 20116 20323
rect 19956 18323 20116 20205
rect 19956 18205 19977 18323
rect 20095 18205 20116 18323
rect 19956 16323 20116 18205
rect 19956 16205 19977 16323
rect 20095 16205 20116 16323
rect 19956 14323 20116 16205
rect 19956 14205 19977 14323
rect 20095 14205 20116 14323
rect 19956 12323 20116 14205
rect 19956 12205 19977 12323
rect 20095 12205 20116 12323
rect 19956 10323 20116 12205
rect 19956 10205 19977 10323
rect 20095 10205 20116 10323
rect 19956 8323 20116 10205
rect 19956 8205 19977 8323
rect 20095 8205 20116 8323
rect 19956 6323 20116 8205
rect 19956 6205 19977 6323
rect 20095 6205 20116 6323
rect 17956 4205 17977 4323
rect 18095 4205 18116 4323
rect 17956 4184 18116 4205
rect 19956 4323 20116 6205
rect 20956 27323 21116 29205
rect 22956 29323 23116 29344
rect 22956 29205 22977 29323
rect 23095 29205 23116 29323
rect 20956 27205 20977 27323
rect 21095 27205 21116 27323
rect 20956 25323 21116 27205
rect 20956 25205 20977 25323
rect 21095 25205 21116 25323
rect 20956 23323 21116 25205
rect 20956 23205 20977 23323
rect 21095 23205 21116 23323
rect 20956 21323 21116 23205
rect 20956 21205 20977 21323
rect 21095 21205 21116 21323
rect 20956 19323 21116 21205
rect 20956 19205 20977 19323
rect 21095 19205 21116 19323
rect 20956 17323 21116 19205
rect 20956 17205 20977 17323
rect 21095 17205 21116 17323
rect 20956 15323 21116 17205
rect 20956 15205 20977 15323
rect 21095 15205 21116 15323
rect 20956 13323 21116 15205
rect 20956 13205 20977 13323
rect 21095 13205 21116 13323
rect 20956 11323 21116 13205
rect 20956 11205 20977 11323
rect 21095 11205 21116 11323
rect 20956 9323 21116 11205
rect 20956 9205 20977 9323
rect 21095 9205 21116 9323
rect 20956 7323 21116 9205
rect 20956 7205 20977 7323
rect 21095 7205 21116 7323
rect 20956 5323 21116 7205
rect 20956 5205 20977 5323
rect 21095 5205 21116 5323
rect 20956 5184 21116 5205
rect 21956 28323 22116 28344
rect 21956 28205 21977 28323
rect 22095 28205 22116 28323
rect 21956 26323 22116 28205
rect 21956 26205 21977 26323
rect 22095 26205 22116 26323
rect 21956 24323 22116 26205
rect 21956 24205 21977 24323
rect 22095 24205 22116 24323
rect 21956 22323 22116 24205
rect 21956 22205 21977 22323
rect 22095 22205 22116 22323
rect 21956 20323 22116 22205
rect 21956 20205 21977 20323
rect 22095 20205 22116 20323
rect 21956 18323 22116 20205
rect 21956 18205 21977 18323
rect 22095 18205 22116 18323
rect 21956 16323 22116 18205
rect 21956 16205 21977 16323
rect 22095 16205 22116 16323
rect 21956 14323 22116 16205
rect 21956 14205 21977 14323
rect 22095 14205 22116 14323
rect 21956 12323 22116 14205
rect 21956 12205 21977 12323
rect 22095 12205 22116 12323
rect 21956 10323 22116 12205
rect 21956 10205 21977 10323
rect 22095 10205 22116 10323
rect 21956 8323 22116 10205
rect 21956 8205 21977 8323
rect 22095 8205 22116 8323
rect 21956 6323 22116 8205
rect 21956 6205 21977 6323
rect 22095 6205 22116 6323
rect 19956 4205 19977 4323
rect 20095 4205 20116 4323
rect 19956 4184 20116 4205
rect 21956 4323 22116 6205
rect 22956 27323 23116 29205
rect 24956 29323 25116 29344
rect 24956 29205 24977 29323
rect 25095 29205 25116 29323
rect 22956 27205 22977 27323
rect 23095 27205 23116 27323
rect 22956 25323 23116 27205
rect 22956 25205 22977 25323
rect 23095 25205 23116 25323
rect 22956 23323 23116 25205
rect 22956 23205 22977 23323
rect 23095 23205 23116 23323
rect 22956 21323 23116 23205
rect 22956 21205 22977 21323
rect 23095 21205 23116 21323
rect 22956 19323 23116 21205
rect 22956 19205 22977 19323
rect 23095 19205 23116 19323
rect 22956 17323 23116 19205
rect 22956 17205 22977 17323
rect 23095 17205 23116 17323
rect 22956 15323 23116 17205
rect 22956 15205 22977 15323
rect 23095 15205 23116 15323
rect 22956 13323 23116 15205
rect 22956 13205 22977 13323
rect 23095 13205 23116 13323
rect 22956 11323 23116 13205
rect 22956 11205 22977 11323
rect 23095 11205 23116 11323
rect 22956 9323 23116 11205
rect 22956 9205 22977 9323
rect 23095 9205 23116 9323
rect 22956 7323 23116 9205
rect 22956 7205 22977 7323
rect 23095 7205 23116 7323
rect 22956 5323 23116 7205
rect 22956 5205 22977 5323
rect 23095 5205 23116 5323
rect 22956 5184 23116 5205
rect 23956 28323 24116 28344
rect 23956 28205 23977 28323
rect 24095 28205 24116 28323
rect 23956 26323 24116 28205
rect 23956 26205 23977 26323
rect 24095 26205 24116 26323
rect 23956 24323 24116 26205
rect 23956 24205 23977 24323
rect 24095 24205 24116 24323
rect 23956 22323 24116 24205
rect 23956 22205 23977 22323
rect 24095 22205 24116 22323
rect 23956 20323 24116 22205
rect 23956 20205 23977 20323
rect 24095 20205 24116 20323
rect 23956 18323 24116 20205
rect 23956 18205 23977 18323
rect 24095 18205 24116 18323
rect 23956 16323 24116 18205
rect 23956 16205 23977 16323
rect 24095 16205 24116 16323
rect 23956 14323 24116 16205
rect 23956 14205 23977 14323
rect 24095 14205 24116 14323
rect 23956 12323 24116 14205
rect 23956 12205 23977 12323
rect 24095 12205 24116 12323
rect 23956 10323 24116 12205
rect 23956 10205 23977 10323
rect 24095 10205 24116 10323
rect 23956 8323 24116 10205
rect 23956 8205 23977 8323
rect 24095 8205 24116 8323
rect 23956 6323 24116 8205
rect 23956 6205 23977 6323
rect 24095 6205 24116 6323
rect 21956 4205 21977 4323
rect 22095 4205 22116 4323
rect 21956 4184 22116 4205
rect 23956 4323 24116 6205
rect 24956 27323 25116 29205
rect 26956 29323 27116 29344
rect 26956 29205 26977 29323
rect 27095 29205 27116 29323
rect 24956 27205 24977 27323
rect 25095 27205 25116 27323
rect 24956 25323 25116 27205
rect 24956 25205 24977 25323
rect 25095 25205 25116 25323
rect 24956 23323 25116 25205
rect 24956 23205 24977 23323
rect 25095 23205 25116 23323
rect 24956 21323 25116 23205
rect 24956 21205 24977 21323
rect 25095 21205 25116 21323
rect 24956 19323 25116 21205
rect 24956 19205 24977 19323
rect 25095 19205 25116 19323
rect 24956 17323 25116 19205
rect 24956 17205 24977 17323
rect 25095 17205 25116 17323
rect 24956 15323 25116 17205
rect 24956 15205 24977 15323
rect 25095 15205 25116 15323
rect 24956 13323 25116 15205
rect 24956 13205 24977 13323
rect 25095 13205 25116 13323
rect 24956 11323 25116 13205
rect 24956 11205 24977 11323
rect 25095 11205 25116 11323
rect 24956 9323 25116 11205
rect 24956 9205 24977 9323
rect 25095 9205 25116 9323
rect 24956 7323 25116 9205
rect 24956 7205 24977 7323
rect 25095 7205 25116 7323
rect 24956 5323 25116 7205
rect 24956 5205 24977 5323
rect 25095 5205 25116 5323
rect 24956 5184 25116 5205
rect 25956 28323 26116 28344
rect 25956 28205 25977 28323
rect 26095 28205 26116 28323
rect 25956 26323 26116 28205
rect 25956 26205 25977 26323
rect 26095 26205 26116 26323
rect 25956 24323 26116 26205
rect 25956 24205 25977 24323
rect 26095 24205 26116 24323
rect 25956 22323 26116 24205
rect 25956 22205 25977 22323
rect 26095 22205 26116 22323
rect 25956 20323 26116 22205
rect 25956 20205 25977 20323
rect 26095 20205 26116 20323
rect 25956 18323 26116 20205
rect 25956 18205 25977 18323
rect 26095 18205 26116 18323
rect 25956 16323 26116 18205
rect 25956 16205 25977 16323
rect 26095 16205 26116 16323
rect 25956 14323 26116 16205
rect 25956 14205 25977 14323
rect 26095 14205 26116 14323
rect 25956 12323 26116 14205
rect 25956 12205 25977 12323
rect 26095 12205 26116 12323
rect 25956 10323 26116 12205
rect 25956 10205 25977 10323
rect 26095 10205 26116 10323
rect 25956 8323 26116 10205
rect 25956 8205 25977 8323
rect 26095 8205 26116 8323
rect 25956 6323 26116 8205
rect 25956 6205 25977 6323
rect 26095 6205 26116 6323
rect 23956 4205 23977 4323
rect 24095 4205 24116 4323
rect 23956 4184 24116 4205
rect 25956 4323 26116 6205
rect 26956 27323 27116 29205
rect 28956 29323 29116 29344
rect 28956 29205 28977 29323
rect 29095 29205 29116 29323
rect 26956 27205 26977 27323
rect 27095 27205 27116 27323
rect 26956 25323 27116 27205
rect 26956 25205 26977 25323
rect 27095 25205 27116 25323
rect 26956 23323 27116 25205
rect 26956 23205 26977 23323
rect 27095 23205 27116 23323
rect 26956 21323 27116 23205
rect 26956 21205 26977 21323
rect 27095 21205 27116 21323
rect 26956 19323 27116 21205
rect 26956 19205 26977 19323
rect 27095 19205 27116 19323
rect 26956 17323 27116 19205
rect 26956 17205 26977 17323
rect 27095 17205 27116 17323
rect 26956 15323 27116 17205
rect 26956 15205 26977 15323
rect 27095 15205 27116 15323
rect 26956 13323 27116 15205
rect 26956 13205 26977 13323
rect 27095 13205 27116 13323
rect 26956 11323 27116 13205
rect 26956 11205 26977 11323
rect 27095 11205 27116 11323
rect 26956 9323 27116 11205
rect 26956 9205 26977 9323
rect 27095 9205 27116 9323
rect 26956 7323 27116 9205
rect 26956 7205 26977 7323
rect 27095 7205 27116 7323
rect 26956 5323 27116 7205
rect 26956 5205 26977 5323
rect 27095 5205 27116 5323
rect 26956 5184 27116 5205
rect 27956 28323 28116 28344
rect 27956 28205 27977 28323
rect 28095 28205 28116 28323
rect 27956 26323 28116 28205
rect 27956 26205 27977 26323
rect 28095 26205 28116 26323
rect 27956 24323 28116 26205
rect 27956 24205 27977 24323
rect 28095 24205 28116 24323
rect 27956 22323 28116 24205
rect 27956 22205 27977 22323
rect 28095 22205 28116 22323
rect 27956 20323 28116 22205
rect 27956 20205 27977 20323
rect 28095 20205 28116 20323
rect 27956 18323 28116 20205
rect 27956 18205 27977 18323
rect 28095 18205 28116 18323
rect 27956 16323 28116 18205
rect 27956 16205 27977 16323
rect 28095 16205 28116 16323
rect 27956 14323 28116 16205
rect 27956 14205 27977 14323
rect 28095 14205 28116 14323
rect 27956 12323 28116 14205
rect 27956 12205 27977 12323
rect 28095 12205 28116 12323
rect 27956 10323 28116 12205
rect 27956 10205 27977 10323
rect 28095 10205 28116 10323
rect 27956 8323 28116 10205
rect 27956 8205 27977 8323
rect 28095 8205 28116 8323
rect 27956 6323 28116 8205
rect 27956 6205 27977 6323
rect 28095 6205 28116 6323
rect 25956 4205 25977 4323
rect 26095 4205 26116 4323
rect 25956 4184 26116 4205
rect 27956 4323 28116 6205
rect 28956 27323 29116 29205
rect 28956 27205 28977 27323
rect 29095 27205 29116 27323
rect 28956 25323 29116 27205
rect 28956 25205 28977 25323
rect 29095 25205 29116 25323
rect 28956 23323 29116 25205
rect 28956 23205 28977 23323
rect 29095 23205 29116 23323
rect 28956 21323 29116 23205
rect 28956 21205 28977 21323
rect 29095 21205 29116 21323
rect 28956 19323 29116 21205
rect 28956 19205 28977 19323
rect 29095 19205 29116 19323
rect 28956 17323 29116 19205
rect 28956 17205 28977 17323
rect 29095 17205 29116 17323
rect 28956 15323 29116 17205
rect 28956 15205 28977 15323
rect 29095 15205 29116 15323
rect 28956 13323 29116 15205
rect 28956 13205 28977 13323
rect 29095 13205 29116 13323
rect 28956 11323 29116 13205
rect 28956 11205 28977 11323
rect 29095 11205 29116 11323
rect 28956 9323 29116 11205
rect 28956 9205 28977 9323
rect 29095 9205 29116 9323
rect 28956 7323 29116 9205
rect 28956 7205 28977 7323
rect 29095 7205 29116 7323
rect 28956 5323 29116 7205
rect 28956 5205 28977 5323
rect 29095 5205 29116 5323
rect 28956 5184 29116 5205
rect 27956 4205 27977 4323
rect 28095 4205 28116 4323
rect 27956 4184 28116 4205
rect 8769 630 8770 662
rect 8769 629 8802 630
<< via4 >>
rect 4977 29205 5095 29323
rect 3977 28205 4095 28323
rect 3977 26205 4095 26323
rect 3977 24205 4095 24323
rect 3977 22205 4095 22323
rect 3977 20205 4095 20323
rect 3977 18205 4095 18323
rect 3977 16205 4095 16323
rect 3977 14205 4095 14323
rect 3977 12205 4095 12323
rect 3977 10205 4095 10323
rect 3977 8205 4095 8323
rect 3977 6205 4095 6323
rect 6977 29205 7095 29323
rect 4977 27205 5095 27323
rect 4977 25205 5095 25323
rect 4977 23205 5095 23323
rect 4977 21205 5095 21323
rect 4977 19205 5095 19323
rect 4977 17205 5095 17323
rect 4977 15205 5095 15323
rect 4977 13205 5095 13323
rect 4977 11205 5095 11323
rect 4977 9205 5095 9323
rect 4977 7205 5095 7323
rect 4977 5205 5095 5323
rect 5977 28205 6095 28323
rect 5977 26205 6095 26323
rect 5977 24205 6095 24323
rect 5977 22205 6095 22323
rect 5977 20205 6095 20323
rect 5977 18205 6095 18323
rect 5977 16205 6095 16323
rect 5977 14205 6095 14323
rect 5977 12205 6095 12323
rect 5977 10205 6095 10323
rect 5977 8205 6095 8323
rect 5977 6205 6095 6323
rect 3977 4205 4095 4323
rect 8977 29205 9095 29323
rect 6977 27205 7095 27323
rect 6977 25205 7095 25323
rect 6977 23205 7095 23323
rect 6977 21205 7095 21323
rect 6977 19205 7095 19323
rect 6977 17205 7095 17323
rect 6977 15205 7095 15323
rect 6977 13205 7095 13323
rect 6977 11205 7095 11323
rect 6977 9205 7095 9323
rect 6977 7205 7095 7323
rect 6977 5205 7095 5323
rect 7977 28205 8095 28323
rect 7977 26205 8095 26323
rect 7977 24205 8095 24323
rect 7977 22205 8095 22323
rect 7977 20205 8095 20323
rect 7977 18205 8095 18323
rect 7977 16205 8095 16323
rect 7977 14205 8095 14323
rect 7977 12205 8095 12323
rect 7977 10205 8095 10323
rect 7977 8205 8095 8323
rect 10977 29205 11095 29323
rect 8977 27205 9095 27323
rect 8977 25205 9095 25323
rect 8977 23205 9095 23323
rect 8977 21205 9095 21323
rect 8977 19205 9095 19323
rect 8977 17205 9095 17323
rect 8977 15205 9095 15323
rect 8977 13205 9095 13323
rect 8977 11205 9095 11323
rect 8977 9205 9095 9323
rect 7977 6205 8095 6323
rect 5977 4205 6095 4323
rect 7977 4205 8095 4323
rect 8977 7205 9095 7323
rect 8977 5205 9095 5323
rect 9977 28205 10095 28323
rect 9977 26205 10095 26323
rect 9977 24205 10095 24323
rect 9977 22205 10095 22323
rect 9977 20205 10095 20323
rect 9977 18205 10095 18323
rect 9977 16205 10095 16323
rect 9977 14205 10095 14323
rect 9977 12205 10095 12323
rect 9977 10205 10095 10323
rect 9977 8205 10095 8323
rect 9977 6205 10095 6323
rect 12977 29205 13095 29323
rect 10977 27205 11095 27323
rect 10977 25205 11095 25323
rect 10977 23205 11095 23323
rect 10977 21205 11095 21323
rect 10977 19205 11095 19323
rect 10977 17205 11095 17323
rect 10977 15205 11095 15323
rect 10977 13205 11095 13323
rect 10977 11205 11095 11323
rect 10977 9205 11095 9323
rect 10977 7205 11095 7323
rect 10977 5205 11095 5323
rect 11977 28205 12095 28323
rect 11977 26205 12095 26323
rect 11977 24205 12095 24323
rect 11977 22205 12095 22323
rect 11977 20205 12095 20323
rect 11977 18205 12095 18323
rect 11977 16205 12095 16323
rect 11977 14205 12095 14323
rect 11977 12205 12095 12323
rect 11977 10205 12095 10323
rect 11977 8205 12095 8323
rect 11977 6205 12095 6323
rect 9977 4205 10095 4323
rect 14977 29205 15095 29323
rect 12977 27205 13095 27323
rect 12977 25205 13095 25323
rect 12977 23205 13095 23323
rect 12977 21205 13095 21323
rect 12977 19205 13095 19323
rect 12977 17205 13095 17323
rect 12977 15205 13095 15323
rect 12977 13205 13095 13323
rect 12977 11205 13095 11323
rect 12977 9205 13095 9323
rect 12977 7205 13095 7323
rect 12977 5205 13095 5323
rect 13977 28205 14095 28323
rect 13977 26205 14095 26323
rect 13977 24205 14095 24323
rect 13977 22205 14095 22323
rect 13977 20205 14095 20323
rect 13977 18205 14095 18323
rect 13977 16205 14095 16323
rect 13977 14205 14095 14323
rect 13977 12205 14095 12323
rect 13977 10205 14095 10323
rect 13977 8205 14095 8323
rect 13977 6205 14095 6323
rect 11977 4205 12095 4323
rect 16977 29205 17095 29323
rect 14977 27205 15095 27323
rect 14977 25205 15095 25323
rect 14977 23205 15095 23323
rect 14977 21205 15095 21323
rect 14977 19205 15095 19323
rect 14977 17205 15095 17323
rect 14977 15205 15095 15323
rect 14977 13205 15095 13323
rect 14977 11205 15095 11323
rect 14977 9205 15095 9323
rect 14977 7205 15095 7323
rect 14977 5205 15095 5323
rect 15977 28205 16095 28323
rect 15977 26205 16095 26323
rect 15977 24205 16095 24323
rect 15977 22205 16095 22323
rect 15977 20205 16095 20323
rect 15977 18205 16095 18323
rect 15977 16205 16095 16323
rect 15977 14205 16095 14323
rect 15977 12205 16095 12323
rect 18977 29205 19095 29323
rect 16977 27205 17095 27323
rect 16977 25205 17095 25323
rect 16977 23205 17095 23323
rect 16977 21205 17095 21323
rect 16977 19205 17095 19323
rect 16977 17205 17095 17323
rect 16977 15205 17095 15323
rect 16977 13205 17095 13323
rect 16977 11205 17095 11323
rect 15977 10205 16095 10323
rect 15977 8205 16095 8323
rect 15977 6205 16095 6323
rect 13977 4205 14095 4323
rect 16977 9205 17095 9323
rect 16977 7205 17095 7323
rect 16977 5205 17095 5323
rect 17977 28205 18095 28323
rect 17977 26205 18095 26323
rect 17977 24205 18095 24323
rect 17977 22205 18095 22323
rect 17977 20205 18095 20323
rect 17977 18205 18095 18323
rect 17977 16205 18095 16323
rect 17977 14205 18095 14323
rect 17977 12205 18095 12323
rect 17977 10205 18095 10323
rect 17977 8205 18095 8323
rect 17977 6205 18095 6323
rect 15977 4205 16095 4323
rect 20977 29205 21095 29323
rect 18977 27205 19095 27323
rect 18977 25205 19095 25323
rect 18977 23205 19095 23323
rect 18977 21205 19095 21323
rect 18977 19205 19095 19323
rect 18977 17205 19095 17323
rect 18977 15205 19095 15323
rect 18977 13205 19095 13323
rect 18977 11205 19095 11323
rect 18977 9205 19095 9323
rect 18977 7205 19095 7323
rect 18977 5205 19095 5323
rect 19977 28205 20095 28323
rect 19977 26205 20095 26323
rect 19977 24205 20095 24323
rect 19977 22205 20095 22323
rect 19977 20205 20095 20323
rect 19977 18205 20095 18323
rect 19977 16205 20095 16323
rect 19977 14205 20095 14323
rect 19977 12205 20095 12323
rect 19977 10205 20095 10323
rect 19977 8205 20095 8323
rect 19977 6205 20095 6323
rect 17977 4205 18095 4323
rect 22977 29205 23095 29323
rect 20977 27205 21095 27323
rect 20977 25205 21095 25323
rect 20977 23205 21095 23323
rect 20977 21205 21095 21323
rect 20977 19205 21095 19323
rect 20977 17205 21095 17323
rect 20977 15205 21095 15323
rect 20977 13205 21095 13323
rect 20977 11205 21095 11323
rect 20977 9205 21095 9323
rect 20977 7205 21095 7323
rect 20977 5205 21095 5323
rect 21977 28205 22095 28323
rect 21977 26205 22095 26323
rect 21977 24205 22095 24323
rect 21977 22205 22095 22323
rect 21977 20205 22095 20323
rect 21977 18205 22095 18323
rect 21977 16205 22095 16323
rect 21977 14205 22095 14323
rect 21977 12205 22095 12323
rect 21977 10205 22095 10323
rect 21977 8205 22095 8323
rect 21977 6205 22095 6323
rect 19977 4205 20095 4323
rect 24977 29205 25095 29323
rect 22977 27205 23095 27323
rect 22977 25205 23095 25323
rect 22977 23205 23095 23323
rect 22977 21205 23095 21323
rect 22977 19205 23095 19323
rect 22977 17205 23095 17323
rect 22977 15205 23095 15323
rect 22977 13205 23095 13323
rect 22977 11205 23095 11323
rect 22977 9205 23095 9323
rect 22977 7205 23095 7323
rect 22977 5205 23095 5323
rect 23977 28205 24095 28323
rect 23977 26205 24095 26323
rect 23977 24205 24095 24323
rect 23977 22205 24095 22323
rect 23977 20205 24095 20323
rect 23977 18205 24095 18323
rect 23977 16205 24095 16323
rect 23977 14205 24095 14323
rect 23977 12205 24095 12323
rect 23977 10205 24095 10323
rect 23977 8205 24095 8323
rect 23977 6205 24095 6323
rect 21977 4205 22095 4323
rect 26977 29205 27095 29323
rect 24977 27205 25095 27323
rect 24977 25205 25095 25323
rect 24977 23205 25095 23323
rect 24977 21205 25095 21323
rect 24977 19205 25095 19323
rect 24977 17205 25095 17323
rect 24977 15205 25095 15323
rect 24977 13205 25095 13323
rect 24977 11205 25095 11323
rect 24977 9205 25095 9323
rect 24977 7205 25095 7323
rect 24977 5205 25095 5323
rect 25977 28205 26095 28323
rect 25977 26205 26095 26323
rect 25977 24205 26095 24323
rect 25977 22205 26095 22323
rect 25977 20205 26095 20323
rect 25977 18205 26095 18323
rect 25977 16205 26095 16323
rect 25977 14205 26095 14323
rect 25977 12205 26095 12323
rect 25977 10205 26095 10323
rect 25977 8205 26095 8323
rect 25977 6205 26095 6323
rect 23977 4205 24095 4323
rect 28977 29205 29095 29323
rect 26977 27205 27095 27323
rect 26977 25205 27095 25323
rect 26977 23205 27095 23323
rect 26977 21205 27095 21323
rect 26977 19205 27095 19323
rect 26977 17205 27095 17323
rect 26977 15205 27095 15323
rect 26977 13205 27095 13323
rect 26977 11205 27095 11323
rect 26977 9205 27095 9323
rect 26977 7205 27095 7323
rect 26977 5205 27095 5323
rect 27977 28205 28095 28323
rect 27977 26205 28095 26323
rect 27977 24205 28095 24323
rect 27977 22205 28095 22323
rect 27977 20205 28095 20323
rect 27977 18205 28095 18323
rect 27977 16205 28095 16323
rect 27977 14205 28095 14323
rect 27977 12205 28095 12323
rect 27977 10205 28095 10323
rect 27977 8205 28095 8323
rect 27977 6205 28095 6323
rect 25977 4205 26095 4323
rect 28977 27205 29095 27323
rect 28977 25205 29095 25323
rect 28977 23205 29095 23323
rect 28977 21205 29095 21323
rect 28977 19205 29095 19323
rect 28977 17205 29095 17323
rect 28977 15205 29095 15323
rect 28977 13205 29095 13323
rect 28977 11205 29095 11323
rect 28977 9205 29095 9323
rect 28977 7205 29095 7323
rect 28977 5205 29095 5323
rect 27977 4205 28095 4323
<< metal5 >>
rect 4956 29323 29116 29344
rect 4956 29205 4977 29323
rect 5095 29205 6977 29323
rect 7095 29205 8977 29323
rect 9095 29205 10977 29323
rect 11095 29205 12977 29323
rect 13095 29205 14977 29323
rect 15095 29205 16977 29323
rect 17095 29205 18977 29323
rect 19095 29205 20977 29323
rect 21095 29205 22977 29323
rect 23095 29205 24977 29323
rect 25095 29205 26977 29323
rect 27095 29205 28977 29323
rect 29095 29205 29116 29323
rect 4956 29184 29116 29205
rect 3956 28323 28116 28344
rect 3956 28205 3977 28323
rect 4095 28205 5977 28323
rect 6095 28205 7977 28323
rect 8095 28205 9977 28323
rect 10095 28205 11977 28323
rect 12095 28205 13977 28323
rect 14095 28205 15977 28323
rect 16095 28205 17977 28323
rect 18095 28205 19977 28323
rect 20095 28205 21977 28323
rect 22095 28205 23977 28323
rect 24095 28205 25977 28323
rect 26095 28205 27977 28323
rect 28095 28205 28116 28323
rect 3956 28184 28116 28205
rect 4956 27323 29116 27344
rect 4956 27205 4977 27323
rect 5095 27205 6977 27323
rect 7095 27205 8977 27323
rect 9095 27205 10977 27323
rect 11095 27205 12977 27323
rect 13095 27205 14977 27323
rect 15095 27205 16977 27323
rect 17095 27205 18977 27323
rect 19095 27205 20977 27323
rect 21095 27205 22977 27323
rect 23095 27205 24977 27323
rect 25095 27205 26977 27323
rect 27095 27205 28977 27323
rect 29095 27205 29116 27323
rect 4956 27184 29116 27205
rect 3956 26323 28116 26344
rect 3956 26205 3977 26323
rect 4095 26205 5977 26323
rect 6095 26205 7977 26323
rect 8095 26205 9977 26323
rect 10095 26205 11977 26323
rect 12095 26205 13977 26323
rect 14095 26205 15977 26323
rect 16095 26205 17977 26323
rect 18095 26205 19977 26323
rect 20095 26205 21977 26323
rect 22095 26205 23977 26323
rect 24095 26205 25977 26323
rect 26095 26205 27977 26323
rect 28095 26205 28116 26323
rect 3956 26184 28116 26205
rect 4956 25323 29116 25344
rect 4956 25205 4977 25323
rect 5095 25205 6977 25323
rect 7095 25205 8977 25323
rect 9095 25205 10977 25323
rect 11095 25205 12977 25323
rect 13095 25205 14977 25323
rect 15095 25205 16977 25323
rect 17095 25205 18977 25323
rect 19095 25205 20977 25323
rect 21095 25205 22977 25323
rect 23095 25205 24977 25323
rect 25095 25205 26977 25323
rect 27095 25205 28977 25323
rect 29095 25205 29116 25323
rect 4956 25184 29116 25205
rect 3956 24323 28116 24344
rect 3956 24205 3977 24323
rect 4095 24205 5977 24323
rect 6095 24205 7977 24323
rect 8095 24205 9977 24323
rect 10095 24205 11977 24323
rect 12095 24205 13977 24323
rect 14095 24205 15977 24323
rect 16095 24205 17977 24323
rect 18095 24205 19977 24323
rect 20095 24205 21977 24323
rect 22095 24205 23977 24323
rect 24095 24205 25977 24323
rect 26095 24205 27977 24323
rect 28095 24205 28116 24323
rect 3956 24184 28116 24205
rect 4956 23323 29116 23344
rect 4956 23205 4977 23323
rect 5095 23205 6977 23323
rect 7095 23205 8977 23323
rect 9095 23205 10977 23323
rect 11095 23205 12977 23323
rect 13095 23205 14977 23323
rect 15095 23205 16977 23323
rect 17095 23205 18977 23323
rect 19095 23205 20977 23323
rect 21095 23205 22977 23323
rect 23095 23205 24977 23323
rect 25095 23205 26977 23323
rect 27095 23205 28977 23323
rect 29095 23205 29116 23323
rect 4956 23184 29116 23205
rect 3956 22323 28116 22344
rect 3956 22205 3977 22323
rect 4095 22205 5977 22323
rect 6095 22205 7977 22323
rect 8095 22205 9977 22323
rect 10095 22205 11977 22323
rect 12095 22205 13977 22323
rect 14095 22205 15977 22323
rect 16095 22205 17977 22323
rect 18095 22205 19977 22323
rect 20095 22205 21977 22323
rect 22095 22205 23977 22323
rect 24095 22205 25977 22323
rect 26095 22205 27977 22323
rect 28095 22205 28116 22323
rect 3956 22184 28116 22205
rect 4956 21323 29116 21344
rect 4956 21205 4977 21323
rect 5095 21205 6977 21323
rect 7095 21205 8977 21323
rect 9095 21205 10977 21323
rect 11095 21205 12977 21323
rect 13095 21205 14977 21323
rect 15095 21205 16977 21323
rect 17095 21205 18977 21323
rect 19095 21205 20977 21323
rect 21095 21205 22977 21323
rect 23095 21205 24977 21323
rect 25095 21205 26977 21323
rect 27095 21205 28977 21323
rect 29095 21205 29116 21323
rect 4956 21184 29116 21205
rect 3956 20323 28116 20344
rect 3956 20205 3977 20323
rect 4095 20205 5977 20323
rect 6095 20205 7977 20323
rect 8095 20205 9977 20323
rect 10095 20205 11977 20323
rect 12095 20205 13977 20323
rect 14095 20205 15977 20323
rect 16095 20205 17977 20323
rect 18095 20205 19977 20323
rect 20095 20205 21977 20323
rect 22095 20205 23977 20323
rect 24095 20205 25977 20323
rect 26095 20205 27977 20323
rect 28095 20205 28116 20323
rect 3956 20184 28116 20205
rect 4956 19323 29116 19344
rect 4956 19205 4977 19323
rect 5095 19205 6977 19323
rect 7095 19205 8977 19323
rect 9095 19205 10977 19323
rect 11095 19205 12977 19323
rect 13095 19205 14977 19323
rect 15095 19205 16977 19323
rect 17095 19205 18977 19323
rect 19095 19205 20977 19323
rect 21095 19205 22977 19323
rect 23095 19205 24977 19323
rect 25095 19205 26977 19323
rect 27095 19205 28977 19323
rect 29095 19205 29116 19323
rect 4956 19184 29116 19205
rect 3956 18323 28116 18344
rect 3956 18205 3977 18323
rect 4095 18205 5977 18323
rect 6095 18205 7977 18323
rect 8095 18205 9977 18323
rect 10095 18205 11977 18323
rect 12095 18205 13977 18323
rect 14095 18205 15977 18323
rect 16095 18205 17977 18323
rect 18095 18205 19977 18323
rect 20095 18205 21977 18323
rect 22095 18205 23977 18323
rect 24095 18205 25977 18323
rect 26095 18205 27977 18323
rect 28095 18205 28116 18323
rect 3956 18184 28116 18205
rect 4956 17323 29116 17344
rect 4956 17205 4977 17323
rect 5095 17205 6977 17323
rect 7095 17205 8977 17323
rect 9095 17205 10977 17323
rect 11095 17205 12977 17323
rect 13095 17205 14977 17323
rect 15095 17205 16977 17323
rect 17095 17205 18977 17323
rect 19095 17205 20977 17323
rect 21095 17205 22977 17323
rect 23095 17205 24977 17323
rect 25095 17205 26977 17323
rect 27095 17205 28977 17323
rect 29095 17205 29116 17323
rect 4956 17184 29116 17205
rect 3956 16323 28116 16344
rect 3956 16205 3977 16323
rect 4095 16205 5977 16323
rect 6095 16205 7977 16323
rect 8095 16205 9977 16323
rect 10095 16205 11977 16323
rect 12095 16205 13977 16323
rect 14095 16205 15977 16323
rect 16095 16205 17977 16323
rect 18095 16205 19977 16323
rect 20095 16205 21977 16323
rect 22095 16205 23977 16323
rect 24095 16205 25977 16323
rect 26095 16205 27977 16323
rect 28095 16205 28116 16323
rect 3956 16184 28116 16205
rect 4956 15323 29116 15344
rect 4956 15205 4977 15323
rect 5095 15205 6977 15323
rect 7095 15205 8977 15323
rect 9095 15205 10977 15323
rect 11095 15205 12977 15323
rect 13095 15205 14977 15323
rect 15095 15205 16977 15323
rect 17095 15205 18977 15323
rect 19095 15205 20977 15323
rect 21095 15205 22977 15323
rect 23095 15205 24977 15323
rect 25095 15205 26977 15323
rect 27095 15205 28977 15323
rect 29095 15205 29116 15323
rect 4956 15184 29116 15205
rect 3956 14323 28116 14344
rect 3956 14205 3977 14323
rect 4095 14205 5977 14323
rect 6095 14205 7977 14323
rect 8095 14205 9977 14323
rect 10095 14205 11977 14323
rect 12095 14205 13977 14323
rect 14095 14205 15977 14323
rect 16095 14205 17977 14323
rect 18095 14205 19977 14323
rect 20095 14205 21977 14323
rect 22095 14205 23977 14323
rect 24095 14205 25977 14323
rect 26095 14205 27977 14323
rect 28095 14205 28116 14323
rect 3956 14184 28116 14205
rect 4956 13323 29116 13344
rect 4956 13205 4977 13323
rect 5095 13205 6977 13323
rect 7095 13205 8977 13323
rect 9095 13205 10977 13323
rect 11095 13205 12977 13323
rect 13095 13205 14977 13323
rect 15095 13205 16977 13323
rect 17095 13205 18977 13323
rect 19095 13205 20977 13323
rect 21095 13205 22977 13323
rect 23095 13205 24977 13323
rect 25095 13205 26977 13323
rect 27095 13205 28977 13323
rect 29095 13205 29116 13323
rect 4956 13184 29116 13205
rect 3956 12323 28116 12344
rect 3956 12205 3977 12323
rect 4095 12205 5977 12323
rect 6095 12205 7977 12323
rect 8095 12205 9977 12323
rect 10095 12205 11977 12323
rect 12095 12205 13977 12323
rect 14095 12205 15977 12323
rect 16095 12205 17977 12323
rect 18095 12205 19977 12323
rect 20095 12205 21977 12323
rect 22095 12205 23977 12323
rect 24095 12205 25977 12323
rect 26095 12205 27977 12323
rect 28095 12205 28116 12323
rect 3956 12184 28116 12205
rect 4956 11323 29116 11344
rect 4956 11205 4977 11323
rect 5095 11205 6977 11323
rect 7095 11205 8977 11323
rect 9095 11205 10977 11323
rect 11095 11205 12977 11323
rect 13095 11205 14977 11323
rect 15095 11205 16977 11323
rect 17095 11205 18977 11323
rect 19095 11205 20977 11323
rect 21095 11205 22977 11323
rect 23095 11205 24977 11323
rect 25095 11205 26977 11323
rect 27095 11205 28977 11323
rect 29095 11205 29116 11323
rect 4956 11184 29116 11205
rect 3956 10323 28116 10344
rect 3956 10205 3977 10323
rect 4095 10205 5977 10323
rect 6095 10205 7977 10323
rect 8095 10205 9977 10323
rect 10095 10205 11977 10323
rect 12095 10205 13977 10323
rect 14095 10205 15977 10323
rect 16095 10205 17977 10323
rect 18095 10205 19977 10323
rect 20095 10205 21977 10323
rect 22095 10205 23977 10323
rect 24095 10205 25977 10323
rect 26095 10205 27977 10323
rect 28095 10205 28116 10323
rect 3956 10184 28116 10205
rect 4956 9323 29116 9344
rect 4956 9205 4977 9323
rect 5095 9205 6977 9323
rect 7095 9205 8977 9323
rect 9095 9205 10977 9323
rect 11095 9205 12977 9323
rect 13095 9205 14977 9323
rect 15095 9205 16977 9323
rect 17095 9205 18977 9323
rect 19095 9205 20977 9323
rect 21095 9205 22977 9323
rect 23095 9205 24977 9323
rect 25095 9205 26977 9323
rect 27095 9205 28977 9323
rect 29095 9205 29116 9323
rect 4956 9184 29116 9205
rect 3956 8323 28116 8344
rect 3956 8205 3977 8323
rect 4095 8205 5977 8323
rect 6095 8205 7977 8323
rect 8095 8205 9977 8323
rect 10095 8205 11977 8323
rect 12095 8205 13977 8323
rect 14095 8205 15977 8323
rect 16095 8205 17977 8323
rect 18095 8205 19977 8323
rect 20095 8205 21977 8323
rect 22095 8205 23977 8323
rect 24095 8205 25977 8323
rect 26095 8205 27977 8323
rect 28095 8205 28116 8323
rect 3956 8184 28116 8205
rect 4956 7323 29116 7344
rect 4956 7205 4977 7323
rect 5095 7205 6977 7323
rect 7095 7205 8977 7323
rect 9095 7205 10977 7323
rect 11095 7205 12977 7323
rect 13095 7205 14977 7323
rect 15095 7205 16977 7323
rect 17095 7205 18977 7323
rect 19095 7205 20977 7323
rect 21095 7205 22977 7323
rect 23095 7205 24977 7323
rect 25095 7205 26977 7323
rect 27095 7205 28977 7323
rect 29095 7205 29116 7323
rect 4956 7184 29116 7205
rect 3956 6323 28116 6344
rect 3956 6205 3977 6323
rect 4095 6205 5977 6323
rect 6095 6205 7977 6323
rect 8095 6205 9977 6323
rect 10095 6205 11977 6323
rect 12095 6205 13977 6323
rect 14095 6205 15977 6323
rect 16095 6205 17977 6323
rect 18095 6205 19977 6323
rect 20095 6205 21977 6323
rect 22095 6205 23977 6323
rect 24095 6205 25977 6323
rect 26095 6205 27977 6323
rect 28095 6205 28116 6323
rect 3956 6184 28116 6205
rect 4956 5323 29116 5344
rect 4956 5205 4977 5323
rect 5095 5205 6977 5323
rect 7095 5205 8977 5323
rect 9095 5205 10977 5323
rect 11095 5205 12977 5323
rect 13095 5205 14977 5323
rect 15095 5205 16977 5323
rect 17095 5205 18977 5323
rect 19095 5205 20977 5323
rect 21095 5205 22977 5323
rect 23095 5205 24977 5323
rect 25095 5205 26977 5323
rect 27095 5205 28977 5323
rect 29095 5205 29116 5323
rect 4956 5184 29116 5205
rect 3956 4323 28116 4344
rect 3956 4205 3977 4323
rect 4095 4205 5977 4323
rect 6095 4205 7977 4323
rect 8095 4205 9977 4323
rect 10095 4205 11977 4323
rect 12095 4205 13977 4323
rect 14095 4205 15977 4323
rect 16095 4205 17977 4323
rect 18095 4205 19977 4323
rect 20095 4205 21977 4323
rect 22095 4205 23977 4323
rect 24095 4205 25977 4323
rect 26095 4205 27977 4323
rect 28095 4205 28116 4323
rect 3956 4184 28116 4205
use sky130_fd_sc_hd__inv_8  _0594_
timestamp 0
transform 1 0 6256 0 -1 28832
box 0 -24 414 296
use sky130_fd_sc_hd__clkinv_1  _0595_
timestamp 0
transform 1 0 9660 0 -1 28288
box 0 -24 138 296
use sky130_fd_sc_hd__inv_1  _0596_
timestamp 0
transform 1 0 19596 0 1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__inv_6  _0597_
timestamp 0
transform 1 0 22448 0 1 22848
box 0 -24 322 296
use sky130_fd_sc_hd__clkinvlp_2  _0598_
timestamp 0
transform 1 0 17296 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__inv_1  _0599_
timestamp 0
transform 1 0 15916 0 -1 29920
box 0 -24 138 296
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 0
transform 1 0 20562 0 1 25568
box 0 -24 138 296
use sky130_fd_sc_hd__clkinv_1  _0601_
timestamp 0
transform 1 0 23966 0 1 24480
box 0 -24 138 296
use sky130_fd_sc_hd__clkinv_1  _0602_
timestamp 0
transform 1 0 24288 0 -1 24480
box 0 -24 138 296
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 0
transform 1 0 21574 0 1 25568
box 0 -24 138 296
use sky130_fd_sc_hd__inv_1  _0604_
timestamp 0
transform 1 0 8096 0 1 4896
box 0 -24 138 296
use sky130_fd_sc_hd__inv_1  _0605_
timestamp 0
transform 1 0 9614 0 -1 7616
box 0 -24 138 296
use sky130_fd_sc_hd__inv_1  _0606_
timestamp 0
transform 1 0 11178 0 1 5984
box 0 -24 138 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _0607_
timestamp 0
transform 1 0 19228 0 1 28288
box 0 -24 506 296
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 0
transform 1 0 20286 0 1 28288
box 0 -24 414 296
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 0
transform 1 0 20378 0 -1 26656
box 0 -24 414 296
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 0
transform 1 0 5014 0 1 10880
box 0 -24 414 296
use sky130_fd_sc_hd__mux2_1  _0611_
timestamp 0
transform 1 0 13662 0 1 10880
box 0 -24 414 296
use sky130_fd_sc_hd__mux2_1  _0612_
timestamp 0
transform 1 0 20332 0 1 27744
box 0 -24 414 296
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 0
transform 1 0 5152 0 1 28288
box 0 -24 414 296
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 0
transform 1 0 5198 0 -1 11968
box 0 -24 414 296
use sky130_fd_sc_hd__mux2_1  _0615_
timestamp 0
transform 1 0 5198 0 -1 28288
box 0 -24 414 296
use sky130_fd_sc_hd__a31oi_1  _0616_
timestamp 0
transform 1 0 7774 0 -1 5440
box 0 -24 230 296
use sky130_fd_sc_hd__nand2b_1  _0617_
timestamp 0
transform 1 0 8924 0 -1 5440
box 0 -24 230 296
use sky130_fd_sc_hd__nor2_1  _0618_
timestamp 0
transform 1 0 8188 0 -1 5440
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_2  _0619_
timestamp 0
transform 1 0 8510 0 1 5440
box 0 -24 230 296
use sky130_fd_sc_hd__nor4_1  _0620_
timestamp 0
transform 1 0 9016 0 1 9792
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0621_
timestamp 0
transform 1 0 9568 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__a221o_1  _0622_
timestamp 0
transform 1 0 9292 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__a21oi_1  _0623_
timestamp 0
transform 1 0 9246 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__nand2_1  _0624_
timestamp 0
transform 1 0 10028 0 -1 5440
box 0 -24 138 296
use sky130_fd_sc_hd__a21oi_1  _0625_
timestamp 0
transform 1 0 10948 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0626_
timestamp 0
transform 1 0 7682 0 -1 5984
box 0 -24 138 296
use sky130_fd_sc_hd__o32ai_1  _0627_
timestamp 0
transform 1 0 7728 0 1 5440
box 0 -24 322 296
use sky130_fd_sc_hd__o21ai_0  _0628_
timestamp 0
transform 1 0 11546 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__xnor2_1  _0629_
timestamp 0
transform 1 0 8050 0 -1 5984
box 0 -24 322 296
use sky130_fd_sc_hd__o21ai_0  _0630_
timestamp 0
transform 1 0 10166 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__a2111oi_0  _0631_
timestamp 0
transform 1 0 8924 0 -1 8704
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_1  _0632_
timestamp 0
transform 1 0 8924 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__nor4_2  _0633_
timestamp 0
transform 1 0 9844 0 -1 5984
box 0 -24 460 296
use sky130_fd_sc_hd__xor2_1  _0634_
timestamp 0
transform 1 0 5750 0 1 8704
box 0 -24 322 296
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 0
transform 1 0 6026 0 -1 18496
box 0 -24 414 296
use sky130_fd_sc_hd__nor3b_2  _0636_
timestamp 0
transform 1 0 15410 0 -1 28288
box 0 -24 460 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _0637_
timestamp 0
transform 1 0 11914 0 1 27744
box 0 -24 506 296
use sky130_fd_sc_hd__nand2_1  _0638_
timestamp 0
transform 1 0 8878 0 -1 29376
box 0 -24 138 296
use sky130_fd_sc_hd__nand3_1  _0639_
timestamp 0
transform 1 0 10304 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__nand4_1  _0640_
timestamp 0
transform 1 0 10488 0 -1 28288
box 0 -24 230 296
use sky130_fd_sc_hd__nor2_2  _0641_
timestamp 0
transform 1 0 17434 0 1 28832
box 0 -24 230 296
use sky130_fd_sc_hd__nor3_2  _0642_
timestamp 0
transform 1 0 17066 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__or3_4  _0643_
timestamp 0
transform 1 0 16606 0 1 28288
box 0 -24 414 296
use sky130_fd_sc_hd__nand2_1  _0644_
timestamp 0
transform 1 0 10396 0 1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__a21oi_1  _0645_
timestamp 0
transform 1 0 10120 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _0646_
timestamp 0
transform 1 0 11684 0 1 28832
box 0 -24 230 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _0647_
timestamp 0
transform 1 0 9246 0 1 27200
box 0 -24 506 296
use sky130_fd_sc_hd__nand2_2  _0648_
timestamp 0
transform 1 0 10258 0 -1 27744
box 0 -24 230 296
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 0
transform 1 0 11592 0 -1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_2  _0650_
timestamp 0
transform 1 0 11730 0 -1 28288
box 0 -24 322 296
use sky130_fd_sc_hd__nor2_4  _0651_
timestamp 0
transform 1 0 11960 0 -1 27744
box 0 -24 414 296
use sky130_fd_sc_hd__xor2_1  _0652_
timestamp 0
transform 1 0 11086 0 1 28832
box 0 -24 322 296
use sky130_fd_sc_hd__a21oi_1  _0653_
timestamp 0
transform 1 0 11684 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0654_
timestamp 0
transform 1 0 12052 0 1 29376
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0655_
timestamp 0
transform 1 0 10258 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0656_
timestamp 0
transform 1 0 10258 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__nor3_1  _0657_
timestamp 0
transform 1 0 8050 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 0
transform 1 0 7728 0 1 25568
box 0 -24 138 296
use sky130_fd_sc_hd__nor4_1  _0659_
timestamp 0
transform 1 0 8970 0 1 25568
box 0 -24 230 296
use sky130_fd_sc_hd__nand3_4  _0660_
timestamp 0
transform 1 0 8142 0 1 25568
box 0 -24 644 296
use sky130_fd_sc_hd__or3b_4  _0661_
timestamp 0
transform 1 0 15686 0 1 28288
box 0 -24 414 296
use sky130_fd_sc_hd__inv_1  _0662_
timestamp 0
transform 1 0 14076 0 1 28832
box 0 -24 138 296
use sky130_fd_sc_hd__a21oi_1  _0663_
timestamp 0
transform 1 0 15686 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__nand2_1  _0664_
timestamp 0
transform 1 0 15686 0 -1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__nor3_2  _0665_
timestamp 0
transform 1 0 15134 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__nand2_4  _0666_
timestamp 0
transform 1 0 14766 0 1 26112
box 0 -24 414 296
use sky130_fd_sc_hd__nand3_1  _0667_
timestamp 0
transform 1 0 17618 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__xor2_1  _0668_
timestamp 0
transform 1 0 15088 0 -1 26656
box 0 -24 322 296
use sky130_fd_sc_hd__nor2_1  _0669_
timestamp 0
transform 1 0 16468 0 1 27200
box 0 -24 138 296
use sky130_fd_sc_hd__a211oi_1  _0670_
timestamp 0
transform 1 0 16330 0 -1 27200
box 0 -24 276 296
use sky130_fd_sc_hd__nand2b_4  _0671_
timestamp 0
transform 1 0 12926 0 1 26112
box 0 -24 506 296
use sky130_fd_sc_hd__nand2b_4  _0672_
timestamp 0
transform 1 0 12926 0 -1 26112
box 0 -24 506 296
use sky130_fd_sc_hd__nand2_1  _0673_
timestamp 0
transform 1 0 13662 0 1 25568
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0674_
timestamp 0
transform 1 0 13616 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__a31oi_1  _0675_
timestamp 0
transform 1 0 13478 0 -1 26656
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0676_
timestamp 0
transform 1 0 13340 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0677_
timestamp 0
transform 1 0 13340 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _0678_
timestamp 0
transform 1 0 18906 0 -1 27744
box 0 -24 230 296
use sky130_fd_sc_hd__nand2_1  _0679_
timestamp 0
transform 1 0 17664 0 1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__and3_4  _0680_
timestamp 0
transform 1 0 18308 0 -1 27744
box 0 -24 414 296
use sky130_fd_sc_hd__nand2_4  _0681_
timestamp 0
transform 1 0 17066 0 -1 25024
box 0 -24 414 296
use sky130_fd_sc_hd__nand3_2  _0682_
timestamp 0
transform 1 0 17664 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__xor2_1  _0683_
timestamp 0
transform 1 0 17204 0 1 25568
box 0 -24 322 296
use sky130_fd_sc_hd__nor2_1  _0684_
timestamp 0
transform 1 0 18216 0 -1 26656
box 0 -24 138 296
use sky130_fd_sc_hd__a211oi_1  _0685_
timestamp 0
transform 1 0 17710 0 1 26112
box 0 -24 276 296
use sky130_fd_sc_hd__nand2b_4  _0686_
timestamp 0
transform 1 0 17618 0 -1 22304
box 0 -24 506 296
use sky130_fd_sc_hd__nand2b_4  _0687_
timestamp 0
transform 1 0 17526 0 1 21760
box 0 -24 506 296
use sky130_fd_sc_hd__nand2_1  _0688_
timestamp 0
transform 1 0 17480 0 1 22848
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0689_
timestamp 0
transform 1 0 17802 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__a31oi_1  _0690_
timestamp 0
transform 1 0 17618 0 1 22304
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0691_
timestamp 0
transform 1 0 18538 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0692_
timestamp 0
transform 1 0 18492 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0693_
timestamp 0
transform 1 0 15778 0 -1 28832
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0694_
timestamp 0
transform 1 0 16100 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__a31oi_1  _0695_
timestamp 0
transform 1 0 16192 0 1 28832
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0696_
timestamp 0
transform 1 0 21206 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0697_
timestamp 0
transform 1 0 21206 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__o21ai_0  _0698_
timestamp 0
transform 1 0 23598 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0699_
timestamp 0
transform 1 0 23920 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0700_
timestamp 0
transform 1 0 23230 0 1 21760
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0701_
timestamp 0
transform 1 0 24196 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0702_
timestamp 0
transform 1 0 22954 0 1 22304
box 0 -24 138 296
use sky130_fd_sc_hd__nor2_1  _0703_
timestamp 0
transform 1 0 22908 0 -1 10880
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0704_
timestamp 0
transform 1 0 23322 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 0
transform 1 0 23138 0 1 10880
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0706_
timestamp 0
transform 1 0 24104 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0707_
timestamp 0
transform 1 0 24472 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0708_
timestamp 0
transform 1 0 22954 0 1 22848
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0709_
timestamp 0
transform 1 0 24150 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0710_
timestamp 0
transform 1 0 23276 0 1 22304
box 0 -24 138 296
use sky130_fd_sc_hd__nor2_1  _0711_
timestamp 0
transform 1 0 23000 0 1 10336
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0712_
timestamp 0
transform 1 0 23966 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0713_
timestamp 0
transform 1 0 23966 0 1 10880
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_2  _0714_
timestamp 0
transform 1 0 20516 0 -1 14144
box 0 -24 230 296
use sky130_fd_sc_hd__nand3_1  _0715_
timestamp 0
transform 1 0 17756 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_2  _0716_
timestamp 0
transform 1 0 17388 0 1 11968
box 0 -24 230 296
use sky130_fd_sc_hd__nand2_4  _0717_
timestamp 0
transform 1 0 17112 0 1 10336
box 0 -24 414 296
use sky130_fd_sc_hd__a21oi_4  _0718_
timestamp 0
transform 1 0 16790 0 1 10880
box 0 -24 598 296
use sky130_fd_sc_hd__nand3_1  _0719_
timestamp 0
transform 1 0 18308 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_4  _0720_
timestamp 0
transform 1 0 17112 0 1 9792
box 0 -24 414 296
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _0721_
timestamp 0
transform 1 0 17066 0 -1 9792
box 0 -24 230 296
use sky130_fd_sc_hd__nor3_1  _0722_
timestamp 0
transform 1 0 19458 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _0723_
timestamp 0
transform 1 0 19458 0 1 14144
box 0 -24 506 296
use sky130_fd_sc_hd__nand2_2  _0724_
timestamp 0
transform 1 0 19412 0 1 11424
box 0 -24 230 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _0725_
timestamp 0
transform 1 0 16284 0 1 12512
box 0 -24 506 296
use sky130_fd_sc_hd__nand2b_4  _0726_
timestamp 0
transform 1 0 16146 0 -1 13056
box 0 -24 506 296
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 0
transform 1 0 18446 0 -1 11424
box 0 -24 138 296
use sky130_fd_sc_hd__a21oi_1  _0728_
timestamp 0
transform 1 0 18446 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__xor2_1  _0729_
timestamp 0
transform 1 0 18446 0 1 11968
box 0 -24 322 296
use sky130_fd_sc_hd__nand2_1  _0730_
timestamp 0
transform 1 0 18630 0 1 11424
box 0 -24 138 296
use sky130_fd_sc_hd__nand2b_1  _0731_
timestamp 0
transform 1 0 18400 0 -1 13600
box 0 -24 230 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _0732_
timestamp 0
transform 1 0 19826 0 -1 14144
box 0 -24 506 296
use sky130_fd_sc_hd__o31ai_1  _0733_
timestamp 0
transform 1 0 18814 0 -1 13600
box 0 -24 276 296
use sky130_fd_sc_hd__nand3_1  _0734_
timestamp 0
transform 1 0 18630 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__xnor2_1  _0735_
timestamp 0
transform 1 0 18170 0 -1 10880
box 0 -24 322 296
use sky130_fd_sc_hd__nand2_1  _0736_
timestamp 0
transform 1 0 18630 0 1 10336
box 0 -24 138 296
use sky130_fd_sc_hd__nor2_2  _0737_
timestamp 0
transform 1 0 17066 0 -1 8704
box 0 -24 230 296
use sky130_fd_sc_hd__and2_4  _0738_
timestamp 0
transform 1 0 17066 0 -1 5984
box 0 -24 322 296
use sky130_fd_sc_hd__nand2_2  _0739_
timestamp 0
transform 1 0 17066 0 -1 6528
box 0 -24 230 296
use sky130_fd_sc_hd__nand2_4  _0740_
timestamp 0
transform 1 0 19780 0 1 5440
box 0 -24 414 296
use sky130_fd_sc_hd__nand3_1  _0741_
timestamp 0
transform 1 0 15962 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0742_
timestamp 0
transform 1 0 16514 0 -1 6528
box 0 -24 138 296
use sky130_fd_sc_hd__a31oi_1  _0743_
timestamp 0
transform 1 0 15916 0 -1 5440
box 0 -24 230 296
use sky130_fd_sc_hd__nor3_1  _0744_
timestamp 0
transform 1 0 15686 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__nand2b_4  _0745_
timestamp 0
transform 1 0 19826 0 -1 4896
box 0 -24 506 296
use sky130_fd_sc_hd__nand2b_4  _0746_
timestamp 0
transform 1 0 19596 0 1 4896
box 0 -24 506 296
use sky130_fd_sc_hd__nand2_1  _0747_
timestamp 0
transform 1 0 18216 0 -1 7616
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0748_
timestamp 0
transform 1 0 18308 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__a31oi_1  _0749_
timestamp 0
transform 1 0 18446 0 1 4896
box 0 -24 230 296
use sky130_fd_sc_hd__a21oi_1  _0750_
timestamp 0
transform 1 0 16422 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0751_
timestamp 0
transform 1 0 17066 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__nor3_2  _0752_
timestamp 0
transform 1 0 16054 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__nand3_2  _0753_
timestamp 0
transform 1 0 14076 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__a21o_1  _0754_
timestamp 0
transform 1 0 14306 0 -1 8160
box 0 -24 276 296
use sky130_fd_sc_hd__nand2_2  _0755_
timestamp 0
transform 1 0 13662 0 1 7616
box 0 -24 230 296
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 0
transform 1 0 13754 0 -1 9248
box 0 -24 138 296
use sky130_fd_sc_hd__a211oi_1  _0757_
timestamp 0
transform 1 0 14352 0 1 8704
box 0 -24 276 296
use sky130_fd_sc_hd__xnor2_1  _0758_
timestamp 0
transform 1 0 14444 0 -1 9248
box 0 -24 322 296
use sky130_fd_sc_hd__o21ai_0  _0759_
timestamp 0
transform 1 0 14950 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0760_
timestamp 0
transform 1 0 14352 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__o21ai_0  _0761_
timestamp 0
transform 1 0 14352 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0762_
timestamp 0
transform 1 0 14766 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__a31oi_1  _0763_
timestamp 0
transform 1 0 14536 0 -1 29376
box 0 -24 230 296
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 0
transform 1 0 13754 0 1 28832
box 0 -24 138 296
use sky130_fd_sc_hd__nand2b_4  _0765_
timestamp 0
transform 1 0 17480 0 -1 21760
box 0 -24 506 296
use sky130_fd_sc_hd__nor2_4  _0766_
timestamp 0
transform 1 0 17894 0 -1 23392
box 0 -24 414 296
use sky130_fd_sc_hd__xor2_1  _0767_
timestamp 0
transform 1 0 17802 0 -1 23936
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 0
transform 1 0 18446 0 1 24480
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _0769_
timestamp 0
transform 1 0 17710 0 -1 26656
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0770_
timestamp 0
transform 1 0 17480 0 -1 24480
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _0771_
timestamp 0
transform 1 0 17112 0 1 25024
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _0772_
timestamp 0
transform 1 0 17802 0 1 26656
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0773_
timestamp 0
transform 1 0 18216 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__nand2_1  _0774_
timestamp 0
transform 1 0 17986 0 -1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0775_
timestamp 0
transform 1 0 18630 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0776_
timestamp 0
transform 1 0 11822 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0777_
timestamp 0
transform 1 0 12190 0 -1 27200
box 0 -24 138 296
use sky130_fd_sc_hd__nand3b_1  _0778_
timestamp 0
transform 1 0 16974 0 1 28832
box 0 -24 276 296
use sky130_fd_sc_hd__nand2_1  _0779_
timestamp 0
transform 1 0 18078 0 -1 28288
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0780_
timestamp 0
transform 1 0 17066 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__nor3_1  _0781_
timestamp 0
transform 1 0 16330 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__inv_1  _0782_
timestamp 0
transform 1 0 16146 0 1 11968
box 0 -24 138 296
use sky130_fd_sc_hd__a21oi_1  _0783_
timestamp 0
transform 1 0 15778 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0784_
timestamp 0
transform 1 0 15686 0 1 12512
box 0 -24 138 296
use sky130_fd_sc_hd__xor2_1  _0785_
timestamp 0
transform 1 0 15686 0 -1 7072
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0786_
timestamp 0
transform 1 0 15226 0 -1 8160
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _0787_
timestamp 0
transform 1 0 15686 0 1 7616
box 0 -24 322 296
use sky130_fd_sc_hd__and4b_4  _0788_
timestamp 0
transform 1 0 20056 0 -1 8160
box 0 -24 506 296
use sky130_fd_sc_hd__xor2_1  _0789_
timestamp 0
transform 1 0 14030 0 1 7072
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0790_
timestamp 0
transform 1 0 15226 0 -1 7616
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _0791_
timestamp 0
transform 1 0 15180 0 -1 9248
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_1  _0792_
timestamp 0
transform 1 0 15732 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__o21ai_0  _0793_
timestamp 0
transform 1 0 17066 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__o311ai_0  _0794_
timestamp 0
transform 1 0 15686 0 1 8704
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0795_
timestamp 0
transform 1 0 18308 0 -1 8160
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0796_
timestamp 0
transform 1 0 18124 0 -1 8704
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0797_
timestamp 0
transform 1 0 16192 0 -1 7072
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0798_
timestamp 0
transform 1 0 17250 0 1 7616
box 0 -24 322 296
use sky130_fd_sc_hd__nor4bb_1  _0799_
timestamp 0
transform 1 0 17066 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__a21oi_1  _0800_
timestamp 0
transform 1 0 17848 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__nor3_1  _0801_
timestamp 0
transform 1 0 17848 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__and4_4  _0802_
timestamp 0
transform 1 0 18998 0 -1 9792
box 0 -24 414 296
use sky130_fd_sc_hd__o21ai_0  _0803_
timestamp 0
transform 1 0 14306 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0804_
timestamp 0
transform 1 0 13708 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__nand3_4  _0805_
timestamp 0
transform 1 0 18354 0 -1 5984
box 0 -24 644 296
use sky130_fd_sc_hd__nor2_4  _0806_
timestamp 0
transform 1 0 19826 0 -1 5984
box 0 -24 414 296
use sky130_fd_sc_hd__o21ai_0  _0807_
timestamp 0
transform 1 0 16836 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__nand3b_1  _0808_
timestamp 0
transform 1 0 18446 0 1 5440
box 0 -24 276 296
use sky130_fd_sc_hd__nor2_4  _0809_
timestamp 0
transform 1 0 18998 0 -1 6528
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_1  _0810_
timestamp 0
transform 1 0 17342 0 -1 5440
box 0 -24 138 296
use sky130_fd_sc_hd__a22oi_1  _0811_
timestamp 0
transform 1 0 17066 0 -1 12512
box 0 -24 276 296
use sky130_fd_sc_hd__a31oi_1  _0812_
timestamp 0
transform 1 0 17664 0 1 14144
box 0 -24 230 296
use sky130_fd_sc_hd__nor2_1  _0813_
timestamp 0
transform 1 0 16974 0 1 11968
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0814_
timestamp 0
transform 1 0 16652 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 0
transform 1 0 16330 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__and4b_4  _0816_
timestamp 0
transform 1 0 22218 0 1 9792
box 0 -24 506 296
use sky130_fd_sc_hd__nor4bb_4  _0817_
timestamp 0
transform 1 0 22586 0 -1 9792
box 0 -24 920 296
use sky130_fd_sc_hd__and4b_4  _0818_
timestamp 0
transform 1 0 18906 0 -1 9248
box 0 -24 506 296
use sky130_fd_sc_hd__nor4b_4  _0819_
timestamp 0
transform 1 0 22034 0 1 8704
box 0 -24 874 296
use sky130_fd_sc_hd__nor4_4  _0820_
timestamp 0
transform 1 0 22218 0 1 7072
box 0 -24 782 296
use sky130_fd_sc_hd__nor4b_2  _0821_
timestamp 0
transform 1 0 22586 0 -1 8704
box 0 -24 552 296
use sky130_fd_sc_hd__nor4bb_4  _0822_
timestamp 0
transform 1 0 22586 0 -1 9248
box 0 -24 920 296
use sky130_fd_sc_hd__nor4bb_4  _0823_
timestamp 0
transform 1 0 22126 0 1 8160
box 0 -24 920 296
use sky130_fd_sc_hd__nor4b_4  _0824_
timestamp 0
transform 1 0 21206 0 -1 8704
box 0 -24 874 296
use sky130_fd_sc_hd__and4b_4  _0825_
timestamp 0
transform 1 0 20700 0 -1 7616
box 0 -24 506 296
use sky130_fd_sc_hd__nor4bb_4  _0826_
timestamp 0
transform 1 0 22080 0 1 7616
box 0 -24 920 296
use sky130_fd_sc_hd__nor4bb_4  _0827_
timestamp 0
transform 1 0 22126 0 1 9248
box 0 -24 920 296
use sky130_fd_sc_hd__nor4b_4  _0828_
timestamp 0
transform 1 0 20746 0 -1 8160
box 0 -24 874 296
use sky130_fd_sc_hd__nor4bb_4  _0829_
timestamp 0
transform 1 0 18860 0 1 9248
box 0 -24 920 296
use sky130_fd_sc_hd__a222oi_1  _0830_
timestamp 0
transform 1 0 29486 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _0831_
timestamp 0
transform 1 0 27140 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _0832_
timestamp 0
transform 1 0 27094 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0833_
timestamp 0
transform 1 0 29486 0 -1 17408
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0834_
timestamp 0
transform 1 0 25622 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0835_
timestamp 0
transform 1 0 29486 0 1 16320
box 0 -24 276 296
use sky130_fd_sc_hd__and4_4  _0836_
timestamp 0
transform 1 0 28612 0 1 16864
box 0 -24 414 296
use sky130_fd_sc_hd__nand3_2  _0837_
timestamp 0
transform 1 0 28704 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__a21oi_1  _0838_
timestamp 0
transform 1 0 23000 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__a22o_1  _0839_
timestamp 0
transform 1 0 26634 0 -1 12512
box 0 -24 322 296
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 0
transform 1 0 29348 0 -1 14688
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _0841_
timestamp 0
transform 1 0 29486 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 0
transform 1 0 29486 0 1 13600
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _0843_
timestamp 0
transform 1 0 27232 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0844_
timestamp 0
transform 1 0 28612 0 1 13600
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0845_
timestamp 0
transform 1 0 25622 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__a221oi_1  _0846_
timestamp 0
transform 1 0 27140 0 -1 12512
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _0847_
timestamp 0
transform 1 0 26772 0 1 13600
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0848_
timestamp 0
transform 1 0 24150 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_4  _0849_
timestamp 0
transform 1 0 20056 0 1 12512
box 0 -24 414 296
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 0
transform 1 0 27186 0 1 5440
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _0851_
timestamp 0
transform 1 0 25346 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__nand2_2  _0852_
timestamp 0
transform 1 0 26726 0 1 5440
box 0 -24 230 296
use sky130_fd_sc_hd__a222oi_1  _0853_
timestamp 0
transform 1 0 25898 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0854_
timestamp 0
transform 1 0 28704 0 -1 8704
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0855_
timestamp 0
transform 1 0 26910 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 0
transform 1 0 29026 0 -1 7072
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _0857_
timestamp 0
transform 1 0 29486 0 1 7616
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _0858_
timestamp 0
transform 1 0 26956 0 1 9248
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_1  _0859_
timestamp 0
transform 1 0 26680 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__nand2_1  _0860_
timestamp 0
transform 1 0 29394 0 -1 11424
box 0 -24 138 296
use sky130_fd_sc_hd__a22oi_1  _0861_
timestamp 0
transform 1 0 29486 0 1 9248
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _0862_
timestamp 0
transform 1 0 28796 0 1 10336
box 0 -24 276 296
use sky130_fd_sc_hd__nand3_1  _0863_
timestamp 0
transform 1 0 29026 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__a22oi_1  _0864_
timestamp 0
transform 1 0 25254 0 1 9248
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0865_
timestamp 0
transform 1 0 26726 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _0866_
timestamp 0
transform 1 0 24242 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__a22o_1  _0867_
timestamp 0
transform 1 0 24426 0 -1 6528
box 0 -24 322 296
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 0
transform 1 0 24748 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__nand4_1  _0869_
timestamp 0
transform 1 0 24702 0 -1 8160
box 0 -24 230 296
use sky130_fd_sc_hd__o21bai_1  _0870_
timestamp 0
transform 1 0 24334 0 -1 11424
box 0 -24 276 296
use sky130_fd_sc_hd__nand4_1  _0871_
timestamp 0
transform 1 0 23874 0 -1 12512
box 0 -24 230 296
use sky130_fd_sc_hd__nand2_1  _0872_
timestamp 0
transform 1 0 18998 0 -1 20128
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _0873_
timestamp 0
transform 1 0 18768 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__nand2_1  _0874_
timestamp 0
transform 1 0 18768 0 -1 17952
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _0875_
timestamp 0
transform 1 0 21942 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0876_
timestamp 0
transform 1 0 20516 0 1 18496
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0877_
timestamp 0
transform 1 0 21298 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__a22o_1  _0878_
timestamp 0
transform 1 0 20286 0 -1 19584
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _0879_
timestamp 0
transform 1 0 20608 0 -1 20128
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _0880_
timestamp 0
transform 1 0 21206 0 1 18496
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0881_
timestamp 0
transform 1 0 21206 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__a222oi_1  _0882_
timestamp 0
transform 1 0 29394 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _0883_
timestamp 0
transform 1 0 26726 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__nand2_1  _0884_
timestamp 0
transform 1 0 26818 0 -1 20672
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _0885_
timestamp 0
transform 1 0 28014 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0886_
timestamp 0
transform 1 0 27370 0 1 18496
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0887_
timestamp 0
transform 1 0 25760 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0888_
timestamp 0
transform 1 0 29486 0 -1 19040
box 0 -24 276 296
use sky130_fd_sc_hd__nand4_1  _0889_
timestamp 0
transform 1 0 27186 0 1 19040
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_2  _0890_
timestamp 0
transform 1 0 25990 0 1 18496
box 0 -24 322 296
use sky130_fd_sc_hd__a222oi_1  _0891_
timestamp 0
transform 1 0 21574 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0892_
timestamp 0
transform 1 0 19964 0 1 15232
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0893_
timestamp 0
transform 1 0 22494 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _0894_
timestamp 0
transform 1 0 22586 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _0895_
timestamp 0
transform 1 0 20102 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0896_
timestamp 0
transform 1 0 22586 0 -1 20672
box 0 -24 276 296
use sky130_fd_sc_hd__and4_4  _0897_
timestamp 0
transform 1 0 22494 0 1 20672
box 0 -24 414 296
use sky130_fd_sc_hd__a31oi_1  _0898_
timestamp 0
transform 1 0 22724 0 1 15232
box 0 -24 230 296
use sky130_fd_sc_hd__a22oi_1  _0899_
timestamp 0
transform 1 0 23966 0 1 16320
box 0 -24 276 296
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 0
transform 1 0 25392 0 -1 22304
box 0 -24 322 296
use sky130_fd_sc_hd__a21oi_1  _0901_
timestamp 0
transform 1 0 25714 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__a22oi_1  _0902_
timestamp 0
transform 1 0 25346 0 -1 19040
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _0903_
timestamp 0
transform 1 0 24564 0 1 20672
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0904_
timestamp 0
transform 1 0 24012 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _0905_
timestamp 0
transform 1 0 24288 0 -1 18496
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _0906_
timestamp 0
transform 1 0 24288 0 -1 20128
box 0 -24 276 296
use sky130_fd_sc_hd__and4_1  _0907_
timestamp 0
transform 1 0 24196 0 -1 19040
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _0908_
timestamp 0
transform 1 0 24702 0 -1 19040
box 0 -24 230 296
use sky130_fd_sc_hd__a21oi_1  _0909_
timestamp 0
transform 1 0 22862 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__nand4_1  _0910_
timestamp 0
transform 1 0 21344 0 -1 14144
box 0 -24 230 296
use sky130_fd_sc_hd__a22oi_1  _0911_
timestamp 0
transform 1 0 22494 0 1 10880
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _0912_
timestamp 0
transform 1 0 21528 0 -1 11968
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0913_
timestamp 0
transform 1 0 22586 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__nand3_1  _0914_
timestamp 0
transform 1 0 21942 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__a222oi_1  _0915_
timestamp 0
transform 1 0 22586 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__a21oi_1  _0916_
timestamp 0
transform 1 0 20194 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__a22oi_1  _0917_
timestamp 0
transform 1 0 20516 0 1 9248
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _0918_
timestamp 0
transform 1 0 22126 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__nand4_1  _0919_
timestamp 0
transform 1 0 20516 0 -1 9792
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0920_
timestamp 0
transform 1 0 19826 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__nand3_1  _0921_
timestamp 0
transform 1 0 19136 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__a31oi_1  _0922_
timestamp 0
transform 1 0 19182 0 -1 13056
box 0 -24 230 296
use sky130_fd_sc_hd__o21ai_0  _0923_
timestamp 0
transform 1 0 15962 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__o21ai_0  _0924_
timestamp 0
transform 1 0 21574 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0925_
timestamp 0
transform 1 0 21298 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__nand2_1  _0926_
timestamp 0
transform 1 0 11592 0 1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 0
transform 1 0 11592 0 1 26112
box 0 -24 138 296
use sky130_fd_sc_hd__nor2_1  _0928_
timestamp 0
transform 1 0 12098 0 1 26112
box 0 -24 138 296
use sky130_fd_sc_hd__nor2_1  _0929_
timestamp 0
transform 1 0 12190 0 1 26656
box 0 -24 138 296
use sky130_fd_sc_hd__a21oi_1  _0930_
timestamp 0
transform 1 0 15686 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0931_
timestamp 0
transform 1 0 15134 0 1 28832
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _0932_
timestamp 0
transform 1 0 18446 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0933_
timestamp 0
transform 1 0 18446 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__xor2_1  _0934_
timestamp 0
transform 1 0 18630 0 -1 25024
box 0 -24 322 296
use sky130_fd_sc_hd__o21ai_0  _0935_
timestamp 0
transform 1 0 18262 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _0936_
timestamp 0
transform 1 0 19090 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__xnor2_1  _0937_
timestamp 0
transform 1 0 10442 0 -1 26656
box 0 -24 322 296
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 0
transform 1 0 10626 0 -1 27200
box 0 -24 230 296
use sky130_fd_sc_hd__nand2b_1  _0939_
timestamp 0
transform 1 0 14858 0 1 26656
box 0 -24 230 296
use sky130_fd_sc_hd__xnor2_1  _0940_
timestamp 0
transform 1 0 18584 0 -1 25568
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0941_
timestamp 0
transform 1 0 16146 0 -1 26656
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _0942_
timestamp 0
transform 1 0 16100 0 1 25568
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_1  _0943_
timestamp 0
transform 1 0 15778 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__or4_1  _0944_
timestamp 0
transform 1 0 16192 0 1 26112
box 0 -24 276 296
use sky130_fd_sc_hd__a21oi_1  _0945_
timestamp 0
transform 1 0 14950 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__nand3b_1  _0946_
timestamp 0
transform 1 0 14812 0 1 25024
box 0 -24 276 296
use sky130_fd_sc_hd__nor2_4  _0947_
timestamp 0
transform 1 0 13386 0 1 22304
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0948_
timestamp 0
transform 1 0 14628 0 -1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nand3b_1  _0949_
timestamp 0
transform 1 0 15778 0 -1 25024
box 0 -24 276 296
use sky130_fd_sc_hd__nor3_4  _0950_
timestamp 0
transform 1 0 15916 0 -1 24480
box 0 -24 598 296
use sky130_fd_sc_hd__nor2_4  _0951_
timestamp 0
transform 1 0 13386 0 -1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 0
transform 1 0 17848 0 1 6528
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_4  _0953_
timestamp 0
transform 1 0 18124 0 -1 6528
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0954_
timestamp 0
transform 1 0 19044 0 1 7616
box 0 -24 414 296
use sky130_fd_sc_hd__or3_4  _0955_
timestamp 0
transform 1 0 17940 0 -1 7072
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0956_
timestamp 0
transform 1 0 20102 0 -1 7616
box 0 -24 414 296
use sky130_fd_sc_hd__or3b_4  _0957_
timestamp 0
transform 1 0 14766 0 1 24480
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0958_
timestamp 0
transform 1 0 14812 0 -1 23936
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0959_
timestamp 0
transform 1 0 18538 0 1 7072
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0960_
timestamp 0
transform 1 0 12972 0 1 23392
box 0 -24 414 296
use sky130_fd_sc_hd__nand3_4  _0961_
timestamp 0
transform 1 0 14812 0 -1 25024
box 0 -24 644 296
use sky130_fd_sc_hd__nor3_4  _0962_
timestamp 0
transform 1 0 13846 0 1 23936
box 0 -24 598 296
use sky130_fd_sc_hd__nor3_4  _0963_
timestamp 0
transform 1 0 13616 0 1 24480
box 0 -24 598 296
use sky130_fd_sc_hd__nor2_4  _0964_
timestamp 0
transform 1 0 12788 0 -1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0965_
timestamp 0
transform 1 0 12972 0 -1 23392
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0966_
timestamp 0
transform 1 0 12834 0 -1 23936
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0967_
timestamp 0
transform 1 0 18860 0 -1 7616
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0968_
timestamp 0
transform 1 0 19872 0 1 7616
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _0969_
timestamp 0
transform 1 0 19596 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _0970_
timestamp 0
transform 1 0 18906 0 1 6528
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _0971_
timestamp 0
transform 1 0 19504 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _0972_
timestamp 0
transform 1 0 21206 0 1 7616
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0973_
timestamp 0
transform 1 0 19918 0 -1 5440
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _0974_
timestamp 0
transform 1 0 20102 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _0975_
timestamp 0
transform 1 0 20194 0 -1 6528
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _0976_
timestamp 0
transform 1 0 19872 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _0977_
timestamp 0
transform 1 0 18998 0 -1 23392
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_4  _0978_
timestamp 0
transform 1 0 12834 0 -1 25024
box 0 -24 598 296
use sky130_fd_sc_hd__nor2_4  _0979_
timestamp 0
transform 1 0 14812 0 1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0980_
timestamp 0
transform 1 0 13018 0 1 24480
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0981_
timestamp 0
transform 1 0 13340 0 1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0982_
timestamp 0
transform 1 0 14582 0 -1 23392
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _0983_
timestamp 0
transform 1 0 19550 0 1 6528
box 0 -24 414 296
use sky130_fd_sc_hd__xor2_1  _0984_
timestamp 0
transform 1 0 19964 0 -1 22848
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _0985_
timestamp 0
transform 1 0 21298 0 -1 25024
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0986_
timestamp 0
transform 1 0 20240 0 1 25024
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0987_
timestamp 0
transform 1 0 20240 0 -1 25024
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_2  _0988_
timestamp 0
transform 1 0 18538 0 1 3808
box 0 -24 598 296
use sky130_fd_sc_hd__xnor2_1  _0989_
timestamp 0
transform 1 0 19090 0 -1 22848
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _0990_
timestamp 0
transform 1 0 19596 0 1 22848
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_2  _0991_
timestamp 0
transform 1 0 20102 0 1 22848
box 0 -24 598 296
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 0
transform 1 0 10396 0 -1 7616
box 0 -24 138 296
use sky130_fd_sc_hd__a21oi_1  _0993_
timestamp 0
transform 1 0 10948 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__o21a_1  _0994_
timestamp 0
transform 1 0 11868 0 1 7072
box 0 -24 276 296
use sky130_fd_sc_hd__a21oi_1  _0995_
timestamp 0
transform 1 0 11546 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__and3_4  _0996_
timestamp 0
transform 1 0 10718 0 -1 7616
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_1  _0997_
timestamp 0
transform 1 0 10718 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _0998_
timestamp 0
transform 1 0 10902 0 -1 8704
box 0 -24 138 296
use sky130_fd_sc_hd__a211oi_1  _0999_
timestamp 0
transform 1 0 10442 0 -1 8704
box 0 -24 276 296
use sky130_fd_sc_hd__a21oi_1  _1000_
timestamp 0
transform 1 0 8188 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__and3_4  _1001_
timestamp 0
transform 1 0 8832 0 1 7072
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_1  _1002_
timestamp 0
transform 1 0 7912 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _1003_
timestamp 0
transform 1 0 6026 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__o21a_1  _1004_
timestamp 0
transform 1 0 6026 0 -1 7072
box 0 -24 276 296
use sky130_fd_sc_hd__a21oi_1  _1005_
timestamp 0
transform 1 0 5934 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__a311oi_1  _1006_
timestamp 0
transform 1 0 6026 0 -1 6528
box 0 -24 322 296
use sky130_fd_sc_hd__and4_4  _1007_
timestamp 0
transform 1 0 7406 0 1 5984
box 0 -24 414 296
use sky130_fd_sc_hd__a31oi_1  _1008_
timestamp 0
transform 1 0 6762 0 1 5984
box 0 -24 230 296
use sky130_fd_sc_hd__nor3_1  _1009_
timestamp 0
transform 1 0 6808 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__o21bai_1  _1010_
timestamp 0
transform 1 0 6394 0 -1 8160
box 0 -24 276 296
use sky130_fd_sc_hd__a21oi_1  _1011_
timestamp 0
transform 1 0 6808 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__a21oi_1  _1012_
timestamp 0
transform 1 0 8096 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__a311oi_1  _1013_
timestamp 0
transform 1 0 7406 0 1 7616
box 0 -24 322 296
use sky130_fd_sc_hd__and4_4  _1014_
timestamp 0
transform 1 0 7636 0 -1 8704
box 0 -24 414 296
use sky130_fd_sc_hd__a31oi_1  _1015_
timestamp 0
transform 1 0 7590 0 1 8704
box 0 -24 230 296
use sky130_fd_sc_hd__nor2_1  _1016_
timestamp 0
transform 1 0 8004 0 1 8704
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_1  _1017_
timestamp 0
transform 1 0 7452 0 1 9792
box 0 -24 138 296
use sky130_fd_sc_hd__xor2_1  _1018_
timestamp 0
transform 1 0 7820 0 -1 9792
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _1019_
timestamp 0
transform 1 0 7958 0 -1 10336
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _1020_
timestamp 0
transform 1 0 8786 0 -1 9792
box 0 -24 230 296
use sky130_fd_sc_hd__a31oi_1  _1021_
timestamp 0
transform 1 0 8326 0 1 10336
box 0 -24 230 296
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _1022_
timestamp 0
transform 1 0 8832 0 -1 10336
box 0 -24 230 296
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _1023_
timestamp 0
transform 1 0 9476 0 -1 9792
box 0 -24 230 296
use sky130_fd_sc_hd__xnor2_1  _1024_
timestamp 0
transform 1 0 9430 0 1 9792
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _1025_
timestamp 0
transform 1 0 9890 0 -1 9792
box 0 -24 322 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _1026_
timestamp 0
transform 1 0 18446 0 -1 15232
box 0 -24 506 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _1027_
timestamp 0
transform 1 0 15732 0 -1 10880
box 0 -24 506 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _1028_
timestamp 0
transform 1 0 11684 0 -1 10880
box 0 -24 506 296
use sky130_fd_sc_hd__nor3_2  _1029_
timestamp 0
transform 1 0 16836 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__nand2_4  _1030_
timestamp 0
transform 1 0 16606 0 1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _1031_
timestamp 0
transform 1 0 15732 0 -1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _1032_
timestamp 0
transform 1 0 16238 0 -1 23392
box 0 -24 414 296
use sky130_fd_sc_hd__nor4_4  _1033_
timestamp 0
transform 1 0 16560 0 1 24480
box 0 -24 782 296
use sky130_fd_sc_hd__nand2b_4  _1034_
timestamp 0
transform 1 0 16376 0 1 21216
box 0 -24 506 296
use sky130_fd_sc_hd__nor2_4  _1035_
timestamp 0
transform 1 0 14904 0 -1 22304
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _1036_
timestamp 0
transform 1 0 16284 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__nor3_2  _1037_
timestamp 0
transform 1 0 16836 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _1038_
timestamp 0
transform 1 0 16146 0 1 22304
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _1039_
timestamp 0
transform 1 0 18170 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _1040_
timestamp 0
transform 1 0 14858 0 1 21760
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _1041_
timestamp 0
transform 1 0 17066 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _1042_
timestamp 0
transform 1 0 15962 0 1 22848
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_4  _1043_
timestamp 0
transform 1 0 14766 0 1 22304
box 0 -24 414 296
use sky130_fd_sc_hd__nor3_2  _1044_
timestamp 0
transform 1 0 16146 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__nor2_4  _1045_
timestamp 0
transform 1 0 14260 0 1 21760
box 0 -24 414 296
use sky130_fd_sc_hd__a222oi_1  _1046_
timestamp 0
transform 1 0 8096 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__a22o_1  _1047_
timestamp 0
transform 1 0 7636 0 -1 20672
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1048_
timestamp 0
transform 1 0 6486 0 -1 21216
box 0 -24 322 296
use sky130_fd_sc_hd__a22oi_1  _1049_
timestamp 0
transform 1 0 4646 0 1 21216
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _1050_
timestamp 0
transform 1 0 4784 0 -1 21216
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1051_
timestamp 0
transform 1 0 4646 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__nand3_1  _1052_
timestamp 0
transform 1 0 4738 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__a221oi_1  _1053_
timestamp 0
transform 1 0 6440 0 1 21760
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_2  _1054_
timestamp 0
transform 1 0 6394 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _1055_
timestamp 0
transform 1 0 8096 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__a22o_1  _1056_
timestamp 0
transform 1 0 7406 0 1 11424
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1057_
timestamp 0
transform 1 0 7406 0 1 11968
box 0 -24 322 296
use sky130_fd_sc_hd__a22oi_1  _1058_
timestamp 0
transform 1 0 4600 0 -1 13600
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _1059_
timestamp 0
transform 1 0 4646 0 1 13056
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1060_
timestamp 0
transform 1 0 4646 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__nand3_1  _1061_
timestamp 0
transform 1 0 5060 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__a221oi_1  _1062_
timestamp 0
transform 1 0 6164 0 -1 13056
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_1  _1063_
timestamp 0
transform 1 0 6486 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__a222oi_1  _1064_
timestamp 0
transform 1 0 4738 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1065_
timestamp 0
transform 1 0 7728 0 1 24480
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1066_
timestamp 0
transform 1 0 6026 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1067_
timestamp 0
transform 1 0 6256 0 -1 23392
box 0 -24 276 296
use sky130_fd_sc_hd__a22o_1  _1068_
timestamp 0
transform 1 0 4646 0 1 25024
box 0 -24 322 296
use sky130_fd_sc_hd__a21oi_1  _1069_
timestamp 0
transform 1 0 6348 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__a222oi_1  _1070_
timestamp 0
transform 1 0 8694 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__and4_1  _1071_
timestamp 0
transform 1 0 6394 0 1 23392
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_1  _1072_
timestamp 0
transform 1 0 4968 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__a22oi_1  _1073_
timestamp 0
transform 1 0 12926 0 1 18496
box 0 -24 276 296
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp 0
transform 1 0 14766 0 -1 20672
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_1  _1075_
timestamp 0
transform 1 0 16468 0 -1 18496
box 0 -24 138 296
use sky130_fd_sc_hd__a22oi_1  _1076_
timestamp 0
transform 1 0 17066 0 -1 18496
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _1077_
timestamp 0
transform 1 0 15594 0 -1 19040
box 0 -24 276 296
use sky130_fd_sc_hd__nand4_1  _1078_
timestamp 0
transform 1 0 15686 0 1 18496
box 0 -24 230 296
use sky130_fd_sc_hd__a222oi_1  _1079_
timestamp 0
transform 1 0 14214 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__a222oi_1  _1080_
timestamp 0
transform 1 0 17250 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__nand4b_1  _1081_
timestamp 0
transform 1 0 15226 0 -1 20672
box 0 -24 322 296
use sky130_fd_sc_hd__a221o_4  _1082_
timestamp 0
transform 1 0 15594 0 -1 21760
box 0 -24 782 296
use sky130_fd_sc_hd__nand2_1  _1083_
timestamp 0
transform 1 0 12236 0 1 16864
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_1  _1084_
timestamp 0
transform 1 0 12328 0 -1 13600
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _1085_
timestamp 0
transform 1 0 11684 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1086_
timestamp 0
transform 1 0 11822 0 1 11968
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _1087_
timestamp 0
transform 1 0 11546 0 -1 12512
box 0 -24 276 296
use sky130_fd_sc_hd__and3_1  _1088_
timestamp 0
transform 1 0 12006 0 -1 12512
box 0 -24 230 296
use sky130_fd_sc_hd__a222oi_1  _1089_
timestamp 0
transform 1 0 11730 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1090_
timestamp 0
transform 1 0 11546 0 -1 16864
box 0 -24 276 296
use sky130_fd_sc_hd__nand2_1  _1091_
timestamp 0
transform 1 0 12006 0 -1 16864
box 0 -24 138 296
use sky130_fd_sc_hd__a221oi_1  _1092_
timestamp 0
transform 1 0 12144 0 1 14144
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _1093_
timestamp 0
transform 1 0 12282 0 -1 13056
box 0 -24 230 296
use sky130_fd_sc_hd__a22o_1  _1094_
timestamp 0
transform 1 0 6762 0 -1 15232
box 0 -24 322 296
use sky130_fd_sc_hd__a22o_1  _1095_
timestamp 0
transform 1 0 6118 0 -1 16320
box 0 -24 322 296
use sky130_fd_sc_hd__a21oi_1  _1096_
timestamp 0
transform 1 0 6624 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__a22o_1  _1097_
timestamp 0
transform 1 0 4830 0 -1 15232
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1098_
timestamp 0
transform 1 0 4738 0 1 14688
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1099_
timestamp 0
transform 1 0 7406 0 1 14688
box 0 -24 322 296
use sky130_fd_sc_hd__a222oi_1  _1100_
timestamp 0
transform 1 0 8786 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__nand4_1  _1101_
timestamp 0
transform 1 0 6348 0 -1 15232
box 0 -24 230 296
use sky130_fd_sc_hd__a221o_1  _1102_
timestamp 0
transform 1 0 6072 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__nand2_1  _1103_
timestamp 0
transform 1 0 9292 0 1 22848
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 0
transform 1 0 11546 0 -1 23392
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _1105_
timestamp 0
transform 1 0 9338 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1106_
timestamp 0
transform 1 0 10074 0 -1 20128
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _1107_
timestamp 0
transform 1 0 10856 0 1 18496
box 0 -24 276 296
use sky130_fd_sc_hd__and3_4  _1108_
timestamp 0
transform 1 0 10212 0 1 19584
box 0 -24 414 296
use sky130_fd_sc_hd__a222oi_1  _1109_
timestamp 0
transform 1 0 10488 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1110_
timestamp 0
transform 1 0 9154 0 -1 24480
box 0 -24 276 296
use sky130_fd_sc_hd__nand2_1  _1111_
timestamp 0
transform 1 0 9430 0 1 23392
box 0 -24 138 296
use sky130_fd_sc_hd__a221oi_1  _1112_
timestamp 0
transform 1 0 10166 0 1 23392
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _1113_
timestamp 0
transform 1 0 10626 0 -1 23392
box 0 -24 230 296
use sky130_fd_sc_hd__a22o_1  _1114_
timestamp 0
transform 1 0 11730 0 -1 20128
box 0 -24 322 296
use sky130_fd_sc_hd__a222oi_1  _1115_
timestamp 0
transform 1 0 12006 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1116_
timestamp 0
transform 1 0 12006 0 -1 23392
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1117_
timestamp 0
transform 1 0 12374 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__a221oi_1  _1118_
timestamp 0
transform 1 0 12236 0 -1 20128
box 0 -24 322 296
use sky130_fd_sc_hd__a22o_1  _1119_
timestamp 0
transform 1 0 10166 0 1 21760
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1120_
timestamp 0
transform 1 0 10580 0 1 21216
box 0 -24 322 296
use sky130_fd_sc_hd__and3_4  _1121_
timestamp 0
transform 1 0 12926 0 -1 21760
box 0 -24 414 296
use sky130_fd_sc_hd__nand3_2  _1122_
timestamp 0
transform 1 0 12144 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1123_
timestamp 0
transform 1 0 4646 0 1 18496
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1124_
timestamp 0
transform 1 0 8786 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__a22o_1  _1125_
timestamp 0
transform 1 0 6670 0 1 17952
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1126_
timestamp 0
transform 1 0 7406 0 1 17952
box 0 -24 322 296
use sky130_fd_sc_hd__a22oi_1  _1127_
timestamp 0
transform 1 0 4646 0 1 17408
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1128_
timestamp 0
transform 1 0 4830 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__nand3_1  _1129_
timestamp 0
transform 1 0 4692 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__a221oi_1  _1130_
timestamp 0
transform 1 0 6348 0 -1 19040
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_1  _1131_
timestamp 0
transform 1 0 6808 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__nand2_1  _1132_
timestamp 0
transform 1 0 9154 0 -1 13600
box 0 -24 138 296
use sky130_fd_sc_hd__a22o_1  _1133_
timestamp 0
transform 1 0 9522 0 -1 16864
box 0 -24 322 296
use sky130_fd_sc_hd__a222oi_1  _1134_
timestamp 0
transform 1 0 10166 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__a22o_1  _1135_
timestamp 0
transform 1 0 8924 0 -1 11968
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1136_
timestamp 0
transform 1 0 9430 0 -1 11968
box 0 -24 322 296
use sky130_fd_sc_hd__a222oi_1  _1137_
timestamp 0
transform 1 0 7866 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__a21oi_1  _1138_
timestamp 0
transform 1 0 10166 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__a22oi_1  _1139_
timestamp 0
transform 1 0 9614 0 -1 14144
box 0 -24 276 296
use sky130_fd_sc_hd__and4_1  _1140_
timestamp 0
transform 1 0 9476 0 -1 13600
box 0 -24 322 296
use sky130_fd_sc_hd__nand3_1  _1141_
timestamp 0
transform 1 0 10166 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__nand2_1  _1142_
timestamp 0
transform 1 0 15134 0 1 16864
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _1143_
timestamp 0
transform 1 0 14444 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1144_
timestamp 0
transform 1 0 15778 0 1 15232
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _1145_
timestamp 0
transform 1 0 16238 0 1 15232
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1146_
timestamp 0
transform 1 0 14306 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1147_
timestamp 0
transform 1 0 14628 0 1 16864
box 0 -24 276 296
use sky130_fd_sc_hd__a222oi_1  _1148_
timestamp 0
transform 1 0 14674 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__and4_1  _1149_
timestamp 0
transform 1 0 14858 0 -1 16864
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _1150_
timestamp 0
transform 1 0 15962 0 1 14688
box 0 -24 230 296
use sky130_fd_sc_hd__nand2_1  _1151_
timestamp 0
transform 1 0 17066 0 1 16864
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_1  _1152_
timestamp 0
transform 1 0 14812 0 1 11968
box 0 -24 138 296
use sky130_fd_sc_hd__a222oi_1  _1153_
timestamp 0
transform 1 0 13386 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1154_
timestamp 0
transform 1 0 14306 0 -1 11968
box 0 -24 276 296
use sky130_fd_sc_hd__a22oi_1  _1155_
timestamp 0
transform 1 0 14214 0 1 11968
box 0 -24 276 296
use sky130_fd_sc_hd__and3_1  _1156_
timestamp 0
transform 1 0 13892 0 1 12512
box 0 -24 230 296
use sky130_fd_sc_hd__a222oi_1  _1157_
timestamp 0
transform 1 0 14536 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__a22oi_1  _1158_
timestamp 0
transform 1 0 17066 0 -1 16864
box 0 -24 276 296
use sky130_fd_sc_hd__nand2_1  _1159_
timestamp 0
transform 1 0 17204 0 1 16320
box 0 -24 138 296
use sky130_fd_sc_hd__a221oi_1  _1160_
timestamp 0
transform 1 0 15226 0 -1 14144
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _1161_
timestamp 0
transform 1 0 14490 0 1 12512
box 0 -24 230 296
use sky130_fd_sc_hd__a21oi_2  _1162_
timestamp 0
transform 1 0 17158 0 1 27744
box 0 -24 322 296
use sky130_fd_sc_hd__o21ai_0  _1163_
timestamp 0
transform 1 0 13340 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__nor2_1  _1164_
timestamp 0
transform 1 0 13294 0 -1 28288
box 0 -24 138 296
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 0
transform 1 0 12788 0 -1 28288
box 0 -24 138 296
use sky130_fd_sc_hd__a221o_1  _1166_
timestamp 0
transform 1 0 14306 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__a21boi_0  _1167_
timestamp 0
transform 1 0 17618 0 -1 28288
box 0 -24 276 296
use sky130_fd_sc_hd__xnor2_1  _1168_
timestamp 0
transform 1 0 22862 0 -1 24480
box 0 -24 322 296
use sky130_fd_sc_hd__xnor2_1  _1169_
timestamp 0
transform 1 0 23092 0 1 23392
box 0 -24 322 296
use sky130_fd_sc_hd__xor2_1  _1170_
timestamp 0
transform 1 0 20240 0 -1 24480
box 0 -24 322 296
use sky130_fd_sc_hd__o22ai_1  _1171_
timestamp 0
transform 1 0 21482 0 -1 26112
box 0 -24 230 296
use sky130_fd_sc_hd__xor2_1  _1172_
timestamp 0
transform 1 0 20378 0 1 23936
box 0 -24 322 296
use sky130_fd_sc_hd__a2bb2oi_1  _1173_
timestamp 0
transform 1 0 23414 0 -1 25568
box 0 -24 322 296
use sky130_fd_sc_hd__o2bb2ai_1  _1174_
timestamp 0
transform 1 0 22816 0 1 25568
box 0 -24 322 296
use sky130_fd_sc_hd__a221oi_1  _1175_
timestamp 0
transform 1 0 23092 0 -1 26112
box 0 -24 322 296
use sky130_fd_sc_hd__nand4_1  _1176_
timestamp 0
transform 1 0 23368 0 -1 24480
box 0 -24 230 296
use sky130_fd_sc_hd__nor4_2  _1177_
timestamp 0
transform 1 0 20746 0 -1 24480
box 0 -24 460 296
use sky130_fd_sc_hd__nor2_1  _1178_
timestamp 0
transform 1 0 17434 0 -1 11424
box 0 -24 138 296
use sky130_fd_sc_hd__o21ai_0  _1179_
timestamp 0
transform 1 0 17066 0 -1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__o22a_1  _1180_
timestamp 0
transform 1 0 16100 0 1 10880
box 0 -24 322 296
use sky130_fd_sc_hd__o21bai_1  _1181_
timestamp 0
transform 1 0 16054 0 -1 11424
box 0 -24 276 296
use sky130_fd_sc_hd__nor2_1  _1182_
timestamp 0
transform 1 0 8786 0 -1 28832
box 0 -24 138 296
use sky130_fd_sc_hd__nor3_1  _1183_
timestamp 0
transform 1 0 6762 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__nor4_2  _1184_
timestamp 0
transform 1 0 6900 0 -1 26656
box 0 -24 460 296
use sky130_fd_sc_hd__mux2_1  _1185_
timestamp 0
transform 1 0 6026 0 -1 26656
box 0 -24 414 296
use sky130_fd_sc_hd__nor2_1  _1186_
timestamp 0
transform 1 0 8418 0 1 28832
box 0 -24 138 296
use sky130_fd_sc_hd__nor2_1  _1187_
timestamp 0
transform 1 0 7406 0 1 28832
box 0 -24 138 296
use sky130_fd_sc_hd__lpflow_isobufsrc_4  _1188_
timestamp 0
transform 1 0 6486 0 1 26656
box 0 -24 506 296
use sky130_fd_sc_hd__a21boi_0  _1189_
timestamp 0
transform 1 0 7130 0 -1 27744
box 0 -24 276 296
use sky130_fd_sc_hd__a31o_1  _1190_
timestamp 0
transform 1 0 7406 0 1 27200
box 0 -24 322 296
use sky130_fd_sc_hd__nor4b_1  _1191_
timestamp 0
transform 1 0 7406 0 1 26656
box 0 -24 322 296
use sky130_fd_sc_hd__mux2_1  _1192_
timestamp 0
transform 1 0 6670 0 -1 26112
box 0 -24 414 296
use sky130_fd_sc_hd__o31ai_1  _1193_
timestamp 0
transform 1 0 8786 0 -1 28288
box 0 -24 276 296
use sky130_fd_sc_hd__nand3_1  _1194_
timestamp 0
transform 1 0 6854 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__o31ai_1  _1195_
timestamp 0
transform 1 0 8096 0 -1 28832
box 0 -24 276 296
use sky130_fd_sc_hd__nand2b_2  _1196_
timestamp 0
transform 1 0 8602 0 1 27200
box 0 -24 322 296
use sky130_fd_sc_hd__nor3_1  _1197_
timestamp 0
transform 1 0 9246 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__mux2_1  _1198_
timestamp 0
transform 1 0 9062 0 -1 26656
box 0 -24 414 296
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _1199_
timestamp 0
transform 1 0 8142 0 -1 27200
box 0 -24 230 296
use sky130_fd_sc_hd__mux2_1  _1200_
timestamp 0
transform 1 0 7774 0 1 26112
box 0 -24 414 296
use sky130_fd_sc_hd__nand2_1  _1201_
timestamp 0
transform 1 0 6440 0 -1 27744
box 0 -24 138 296
use sky130_fd_sc_hd__lpflow_isobufsrc_1  _1202_
timestamp 0
transform 1 0 6670 0 1 28288
box 0 -24 230 296
use sky130_fd_sc_hd__nor3b_1  _1203_
timestamp 0
transform 1 0 8786 0 -1 27200
box 0 -24 276 296
use sky130_fd_sc_hd__mux2_1  _1204_
timestamp 0
transform 1 0 8326 0 1 26656
box 0 -24 414 296
use sky130_fd_sc_hd__o31ai_1  _1205_
timestamp 0
transform 1 0 8740 0 1 28832
box 0 -24 276 296
use sky130_fd_sc_hd__o31ai_1  _1206_
timestamp 0
transform 1 0 6716 0 1 28832
box 0 -24 276 296
use sky130_fd_sc_hd__mux2_1  _1207_
timestamp 0
transform 1 0 6026 0 -1 27200
box 0 -24 414 296
use sky130_fd_sc_hd__edfxtp_1  _1208_
timestamp 0
transform 1 0 5520 0 1 26112
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1209_
timestamp 0
transform 1 0 6716 0 -1 27200
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1210_
timestamp 0
transform 1 0 6486 0 -1 25568
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1211_
timestamp 0
transform 1 0 8418 0 1 28288
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1212_
timestamp 0
transform 1 0 9062 0 -1 26112
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1213_
timestamp 0
transform 1 0 7268 0 -1 26112
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1214_
timestamp 0
transform 1 0 8418 0 1 26112
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1215_
timestamp 0
transform 1 0 6808 0 -1 29376
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1216_
timestamp 0
transform 1 0 5336 0 1 27200
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1217_
timestamp 0
transform 1 0 4508 0 -1 27200
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1218_
timestamp 0
transform 1 0 4508 0 -1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1219_
timestamp 0
transform 1 0 4508 0 -1 27744
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1220_
timestamp 0
transform 1 0 19136 0 1 27200
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1221_
timestamp 0
transform 1 0 12374 0 -1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1222_
timestamp 0
transform 1 0 4508 0 -1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1223_
timestamp 0
transform 1 0 19136 0 1 26656
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1224_
timestamp 0
transform 1 0 19090 0 1 26112
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1225_
timestamp 0
transform 1 0 5244 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1226_
timestamp 0
transform 1 0 10028 0 -1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1227_
timestamp 0
transform 1 0 16928 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1228_
timestamp 0
transform 1 0 14444 0 -1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__dfrtp_4  _1229_
timestamp 0
transform 1 0 10626 0 1 7072
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1230_
timestamp 0
transform 1 0 10810 0 1 6528
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1231_
timestamp 0
transform 1 0 10534 0 1 7616
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1232_
timestamp 0
transform 1 0 10350 0 1 8704
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1233_
timestamp 0
transform 1 0 7590 0 1 7072
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1234_
timestamp 0
transform 1 0 5520 0 1 7072
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1235_
timestamp 0
transform 1 0 5474 0 1 5984
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1236_
timestamp 0
transform 1 0 6578 0 -1 6528
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1237_
timestamp 0
transform 1 0 6394 0 -1 8704
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1238_
timestamp 0
transform 1 0 6854 0 -1 8160
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 0
transform 1 0 7636 0 1 8160
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_4  _1240_
timestamp 0
transform 1 0 7636 0 1 9248
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1241_
timestamp 0
transform 1 0 7774 0 1 9792
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_1  _1242_
timestamp 0
transform 1 0 8740 0 1 10336
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_4  _1243_
timestamp 0
transform 1 0 9522 0 -1 10336
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 0
transform 1 0 10166 0 1 9792
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_4  _1245_
timestamp 0
transform 1 0 15594 0 -1 10336
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1246_
timestamp 0
transform 1 0 15870 0 1 10336
box 0 -24 1058 296
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 0
transform 1 0 15594 0 -1 12512
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 0
transform 1 0 15916 0 -1 9248
box 0 -24 736 296
use sky130_fd_sc_hd__edfxtp_1  _1249_
timestamp 0
transform 1 0 28106 0 -1 8160
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1250_
timestamp 0
transform 1 0 26726 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1251_
timestamp 0
transform 1 0 28106 0 -1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1252_
timestamp 0
transform 1 0 28106 0 -1 9248
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1253_
timestamp 0
transform 1 0 25806 0 -1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1254_
timestamp 0
transform 1 0 23506 0 -1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1255_
timestamp 0
transform 1 0 17710 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1256_
timestamp 0
transform 1 0 18308 0 -1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1257_
timestamp 0
transform 1 0 19366 0 1 10336
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1258_
timestamp 0
transform 1 0 26726 0 1 8704
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1259_
timestamp 0
transform 1 0 28198 0 -1 22848
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1260_
timestamp 0
transform 1 0 24610 0 1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1261_
timestamp 0
transform 1 0 28106 0 -1 10336
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1262_
timestamp 0
transform 1 0 27968 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1263_
timestamp 0
transform 1 0 24610 0 1 22848
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1264_
timestamp 0
transform 1 0 21206 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1265_
timestamp 0
transform 1 0 21298 0 1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1266_
timestamp 0
transform 1 0 19688 0 1 8704
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1267_
timestamp 0
transform 1 0 25346 0 -1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1268_
timestamp 0
transform 1 0 28198 0 -1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1269_
timestamp 0
transform 1 0 25208 0 1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1270_
timestamp 0
transform 1 0 27508 0 1 10336
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1271_
timestamp 0
transform 1 0 27968 0 1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1272_
timestamp 0
transform 1 0 23138 0 -1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1273_
timestamp 0
transform 1 0 19504 0 1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1274_
timestamp 0
transform 1 0 19320 0 1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1275_
timestamp 0
transform 1 0 21068 0 -1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1276_
timestamp 0
transform 1 0 24058 0 1 4352
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1277_
timestamp 0
transform 1 0 25898 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1278_
timestamp 0
transform 1 0 25852 0 -1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1279_
timestamp 0
transform 1 0 25668 0 -1 7072
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1280_
timestamp 0
transform 1 0 25530 0 -1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1281_
timestamp 0
transform 1 0 22954 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1282_
timestamp 0
transform 1 0 19366 0 1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1283_
timestamp 0
transform 1 0 21206 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1284_
timestamp 0
transform 1 0 21068 0 -1 4896
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1285_
timestamp 0
transform 1 0 27968 0 1 6528
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1286_
timestamp 0
transform 1 0 28290 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1287_
timestamp 0
transform 1 0 25898 0 -1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1288_
timestamp 0
transform 1 0 27968 0 1 9248
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1289_
timestamp 0
transform 1 0 24518 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1290_
timestamp 0
transform 1 0 22448 0 1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1291_
timestamp 0
transform 1 0 17756 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1292_
timestamp 0
transform 1 0 20056 0 -1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1293_
timestamp 0
transform 1 0 21068 0 -1 5440
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1294_
timestamp 0
transform 1 0 25622 0 -1 9248
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1295_
timestamp 0
transform 1 0 24242 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1296_
timestamp 0
transform 1 0 27692 0 1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1297_
timestamp 0
transform 1 0 28106 0 -1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1298_
timestamp 0
transform 1 0 28198 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1299_
timestamp 0
transform 1 0 22724 0 -1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1300_
timestamp 0
transform 1 0 18906 0 1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1301_
timestamp 0
transform 1 0 18308 0 -1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1302_
timestamp 0
transform 1 0 20792 0 -1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1303_
timestamp 0
transform 1 0 28106 0 -1 7616
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1304_
timestamp 0
transform 1 0 27968 0 1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1305_
timestamp 0
transform 1 0 27830 0 1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1306_
timestamp 0
transform 1 0 23966 0 1 9248
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1307_
timestamp 0
transform 1 0 26174 0 -1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1308_
timestamp 0
transform 1 0 24426 0 1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1309_
timestamp 0
transform 1 0 19228 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1310_
timestamp 0
transform 1 0 21206 0 1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1311_
timestamp 0
transform 1 0 19826 0 -1 9248
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1312_
timestamp 0
transform 1 0 27922 0 1 7616
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1313_
timestamp 0
transform 1 0 28198 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1314_
timestamp 0
transform 1 0 28106 0 -1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1315_
timestamp 0
transform 1 0 23966 0 1 6528
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1316_
timestamp 0
transform 1 0 27968 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1317_
timestamp 0
transform 1 0 23000 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1318_
timestamp 0
transform 1 0 18308 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1319_
timestamp 0
transform 1 0 18446 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1320_
timestamp 0
transform 1 0 21068 0 -1 7072
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1321_
timestamp 0
transform 1 0 23782 0 -1 5440
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1322_
timestamp 0
transform 1 0 24334 0 1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1323_
timestamp 0
transform 1 0 24334 0 1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1324_
timestamp 0
transform 1 0 23138 0 -1 6528
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1325_
timestamp 0
transform 1 0 24472 0 1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1326_
timestamp 0
transform 1 0 22816 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1327_
timestamp 0
transform 1 0 20010 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1328_
timestamp 0
transform 1 0 20516 0 -1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1329_
timestamp 0
transform 1 0 20194 0 -1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1330_
timestamp 0
transform 1 0 24610 0 1 10336
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1331_
timestamp 0
transform 1 0 25346 0 -1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1332_
timestamp 0
transform 1 0 24472 0 1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1333_
timestamp 0
transform 1 0 23276 0 -1 7072
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1334_
timestamp 0
transform 1 0 25346 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1335_
timestamp 0
transform 1 0 22954 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1336_
timestamp 0
transform 1 0 20240 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1337_
timestamp 0
transform 1 0 20746 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1338_
timestamp 0
transform 1 0 21206 0 1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1339_
timestamp 0
transform 1 0 28198 0 -1 6528
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1340_
timestamp 0
transform 1 0 28244 0 -1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1341_
timestamp 0
transform 1 0 28336 0 -1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1342_
timestamp 0
transform 1 0 23184 0 -1 8160
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1343_
timestamp 0
transform 1 0 28106 0 -1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1344_
timestamp 0
transform 1 0 22908 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1345_
timestamp 0
transform 1 0 19504 0 1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1346_
timestamp 0
transform 1 0 21068 0 -1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1347_
timestamp 0
transform 1 0 21068 0 -1 6528
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1348_
timestamp 0
transform 1 0 25806 0 -1 8704
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1349_
timestamp 0
transform 1 0 26220 0 -1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1350_
timestamp 0
transform 1 0 26174 0 -1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1351_
timestamp 0
transform 1 0 23828 0 -1 9248
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1352_
timestamp 0
transform 1 0 26266 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1353_
timestamp 0
transform 1 0 24242 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1354_
timestamp 0
transform 1 0 20746 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1355_
timestamp 0
transform 1 0 21068 0 -1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1356_
timestamp 0
transform 1 0 21206 0 1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1357_
timestamp 0
transform 1 0 23966 0 1 4896
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1358_
timestamp 0
transform 1 0 26726 0 1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1359_
timestamp 0
transform 1 0 25990 0 -1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1360_
timestamp 0
transform 1 0 25806 0 -1 7616
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1361_
timestamp 0
transform 1 0 26128 0 -1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1362_
timestamp 0
transform 1 0 23414 0 -1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1363_
timestamp 0
transform 1 0 17710 0 -1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1364_
timestamp 0
transform 1 0 18998 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1365_
timestamp 0
transform 1 0 21206 0 1 4896
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1366_
timestamp 0
transform 1 0 25346 0 -1 10336
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1367_
timestamp 0
transform 1 0 25990 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1368_
timestamp 0
transform 1 0 25346 0 -1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1369_
timestamp 0
transform 1 0 23368 0 -1 8704
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1370_
timestamp 0
transform 1 0 25576 0 -1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1371_
timestamp 0
transform 1 0 23000 0 -1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1372_
timestamp 0
transform 1 0 21206 0 1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1373_
timestamp 0
transform 1 0 21298 0 1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1374_
timestamp 0
transform 1 0 21206 0 1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1375_
timestamp 0
transform 1 0 26404 0 -1 5984
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1376_
timestamp 0
transform 1 0 26726 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1377_
timestamp 0
transform 1 0 25944 0 -1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1378_
timestamp 0
transform 1 0 26726 0 1 7072
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1379_
timestamp 0
transform 1 0 26726 0 1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1380_
timestamp 0
transform 1 0 24380 0 1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1381_
timestamp 0
transform 1 0 21068 0 -1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1382_
timestamp 0
transform 1 0 21068 0 -1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1383_
timestamp 0
transform 1 0 21206 0 1 6528
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1384_
timestamp 0
transform 1 0 19366 0 1 23392
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1385_
timestamp 0
transform 1 0 19550 0 1 24480
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1386_
timestamp 0
transform 1 0 21942 0 1 24480
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1387_
timestamp 0
transform 1 0 21804 0 1 23392
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1388_
timestamp 0
transform 1 0 21712 0 1 23936
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1389_
timestamp 0
transform 1 0 21666 0 1 25024
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1390_
timestamp 0
transform 1 0 20194 0 -1 26112
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1391_
timestamp 0
transform 1 0 21068 0 -1 26656
box 0 -24 1104 296
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 0
transform 1 0 18446 0 1 9792
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 0
transform 1 0 14306 0 -1 10336
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 0
transform 1 0 14030 0 1 9248
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 0
transform 1 0 13432 0 1 8704
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 0
transform 1 0 13708 0 1 6528
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 0
transform 1 0 16560 0 1 4352
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 0
transform 1 0 18400 0 -1 4896
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 0
transform 1 0 14996 0 -1 5440
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 0
transform 1 0 17250 0 1 5440
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 0
transform 1 0 18676 0 -1 10880
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 0
transform 1 0 18676 0 1 13600
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 0
transform 1 0 18676 0 -1 11968
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 0
transform 1 0 17066 0 -1 14144
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 0
transform 1 0 15594 0 -1 13600
box 0 -24 736 296
use sky130_fd_sc_hd__edfxtp_1  _1406_
timestamp 0
transform 1 0 3404 0 -1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1407_
timestamp 0
transform 1 0 3312 0 -1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1408_
timestamp 0
transform 1 0 3358 0 -1 25568
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1409_
timestamp 0
transform 1 0 14168 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1410_
timestamp 0
transform 1 0 10672 0 1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1411_
timestamp 0
transform 1 0 3128 0 1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1412_
timestamp 0
transform 1 0 9016 0 -1 23936
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1413_
timestamp 0
transform 1 0 11086 0 1 24480
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1414_
timestamp 0
transform 1 0 3312 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1415_
timestamp 0
transform 1 0 8464 0 1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1416_
timestamp 0
transform 1 0 13800 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1417_
timestamp 0
transform 1 0 14306 0 -1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 0
transform 1 0 24150 0 -1 10880
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 0
transform 1 0 23230 0 -1 22848
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 0
transform 1 0 24288 0 1 23392
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 0
transform 1 0 23230 0 -1 10880
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 0
transform 1 0 23276 0 -1 22304
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1423_
timestamp 0
transform 1 0 23966 0 -1 23936
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1424_
timestamp 0
transform 1 0 20424 0 -1 23392
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1425_
timestamp 0
transform 1 0 21344 0 -1 23392
box 0 -24 736 296
use sky130_fd_sc_hd__dfrtp_4  _1426_
timestamp 0
transform 1 0 5704 0 1 8160
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1427_
timestamp 0
transform 1 0 12926 0 1 28288
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1428_
timestamp 0
transform 1 0 14214 0 1 28288
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1429_
timestamp 0
transform 1 0 17434 0 -1 28832
box 0 -24 1058 296
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 0
transform 1 0 15916 0 -1 29376
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 0
transform 1 0 14996 0 -1 29376
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 0
transform 1 0 18446 0 1 22304
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 0
transform 1 0 17618 0 -1 22848
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 0
transform 1 0 17802 0 -1 26112
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 0
transform 1 0 18308 0 -1 23936
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 0
transform 1 0 13110 0 1 27200
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 0
transform 1 0 13616 0 1 26112
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 0
transform 1 0 16468 0 1 26656
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 0
transform 1 0 18492 0 1 25024
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 0
transform 1 0 9982 0 -1 29376
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 0
transform 1 0 11638 0 -1 29376
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 0
transform 1 0 10166 0 1 28288
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 0
transform 1 0 10258 0 1 26656
box 0 -24 736 296
use sky130_fd_sc_hd__edfxtp_1  _1444_
timestamp 0
transform 1 0 5520 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1445_
timestamp 0
transform 1 0 5796 0 1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1446_
timestamp 0
transform 1 0 5474 0 1 22848
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1447_
timestamp 0
transform 1 0 15548 0 -1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1448_
timestamp 0
transform 1 0 9936 0 -1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1449_
timestamp 0
transform 1 0 5566 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1450_
timestamp 0
transform 1 0 9982 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1451_
timestamp 0
transform 1 0 11316 0 1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1452_
timestamp 0
transform 1 0 5612 0 1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1453_
timestamp 0
transform 1 0 7268 0 -1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1454_
timestamp 0
transform 1 0 15364 0 -1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1455_
timestamp 0
transform 1 0 12926 0 1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 0
transform 1 0 14582 0 -1 27200
box 0 -24 736 296
use sky130_fd_sc_hd__edfxtp_1  _1457_
timestamp 0
transform 1 0 3772 0 -1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1458_
timestamp 0
transform 1 0 3634 0 -1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1459_
timestamp 0
transform 1 0 4416 0 -1 26112
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1460_
timestamp 0
transform 1 0 11822 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1461_
timestamp 0
transform 1 0 10856 0 1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1462_
timestamp 0
transform 1 0 3772 0 -1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1463_
timestamp 0
transform 1 0 9660 0 -1 25568
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1464_
timestamp 0
transform 1 0 11546 0 -1 25024
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1465_
timestamp 0
transform 1 0 3588 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1466_
timestamp 0
transform 1 0 6946 0 -1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1467_
timestamp 0
transform 1 0 12788 0 -1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1468_
timestamp 0
transform 1 0 12788 0 -1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1469_
timestamp 0
transform 1 0 5152 0 1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1470_
timestamp 0
transform 1 0 5198 0 1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1471_
timestamp 0
transform 1 0 5106 0 1 23392
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1472_
timestamp 0
transform 1 0 14168 0 1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1473_
timestamp 0
transform 1 0 11408 0 1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1474_
timestamp 0
transform 1 0 4508 0 -1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1475_
timestamp 0
transform 1 0 10028 0 -1 22848
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1476_
timestamp 0
transform 1 0 9522 0 -1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1477_
timestamp 0
transform 1 0 5382 0 1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1478_
timestamp 0
transform 1 0 8096 0 1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1479_
timestamp 0
transform 1 0 14168 0 1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1480_
timestamp 0
transform 1 0 12788 0 -1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1481_
timestamp 0
transform 1 0 3128 0 1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1482_
timestamp 0
transform 1 0 3128 0 1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1483_
timestamp 0
transform 1 0 3128 0 1 23936
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1484_
timestamp 0
transform 1 0 16146 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1485_
timestamp 0
transform 1 0 10948 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1486_
timestamp 0
transform 1 0 5704 0 1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1487_
timestamp 0
transform 1 0 8142 0 1 23392
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1488_
timestamp 0
transform 1 0 8648 0 1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1489_
timestamp 0
transform 1 0 3128 0 1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1490_
timestamp 0
transform 1 0 8786 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1491_
timestamp 0
transform 1 0 14674 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1492_
timestamp 0
transform 1 0 15916 0 1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1493_
timestamp 0
transform 1 0 3128 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1494_
timestamp 0
transform 1 0 3128 0 1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1495_
timestamp 0
transform 1 0 6900 0 -1 23936
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1496_
timestamp 0
transform 1 0 14306 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1497_
timestamp 0
transform 1 0 10028 0 -1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1498_
timestamp 0
transform 1 0 3128 0 1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1499_
timestamp 0
transform 1 0 9614 0 -1 25024
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1500_
timestamp 0
transform 1 0 10994 0 1 23392
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1501_
timestamp 0
transform 1 0 3128 0 1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1502_
timestamp 0
transform 1 0 6900 0 -1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1503_
timestamp 0
transform 1 0 13386 0 1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1504_
timestamp 0
transform 1 0 13248 0 1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1505_
timestamp 0
transform 1 0 7590 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1506_
timestamp 0
transform 1 0 7268 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1507_
timestamp 0
transform 1 0 7268 0 -1 22848
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1508_
timestamp 0
transform 1 0 13478 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1509_
timestamp 0
transform 1 0 10856 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1510_
timestamp 0
transform 1 0 7820 0 1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1511_
timestamp 0
transform 1 0 8418 0 1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1512_
timestamp 0
transform 1 0 11408 0 1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1513_
timestamp 0
transform 1 0 7268 0 -1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1514_
timestamp 0
transform 1 0 9200 0 -1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1515_
timestamp 0
transform 1 0 12788 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1516_
timestamp 0
transform 1 0 12466 0 -1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1517_
timestamp 0
transform 1 0 3496 0 -1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1518_
timestamp 0
transform 1 0 5612 0 1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1519_
timestamp 0
transform 1 0 3128 0 1 25024
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1520_
timestamp 0
transform 1 0 11408 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1521_
timestamp 0
transform 1 0 10166 0 1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1522_
timestamp 0
transform 1 0 3542 0 -1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1523_
timestamp 0
transform 1 0 8648 0 1 25024
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1524_
timestamp 0
transform 1 0 10994 0 1 25024
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1525_
timestamp 0
transform 1 0 3128 0 1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1526_
timestamp 0
transform 1 0 6854 0 -1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1527_
timestamp 0
transform 1 0 12604 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1528_
timestamp 0
transform 1 0 12558 0 -1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1529_
timestamp 0
transform 1 0 5336 0 1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1530_
timestamp 0
transform 1 0 3128 0 1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1531_
timestamp 0
transform 1 0 3450 0 -1 24480
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1532_
timestamp 0
transform 1 0 15962 0 1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1533_
timestamp 0
transform 1 0 10028 0 -1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1534_
timestamp 0
transform 1 0 7268 0 -1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1535_
timestamp 0
transform 1 0 10166 0 1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1536_
timestamp 0
transform 1 0 11408 0 1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1537_
timestamp 0
transform 1 0 5474 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1538_
timestamp 0
transform 1 0 8786 0 -1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1539_
timestamp 0
transform 1 0 15318 0 -1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1540_
timestamp 0
transform 1 0 14306 0 -1 12512
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1541_
timestamp 0
transform 1 0 5290 0 1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1542_
timestamp 0
transform 1 0 5336 0 1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1543_
timestamp 0
transform 1 0 5290 0 1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1544_
timestamp 0
transform 1 0 14306 0 -1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1545_
timestamp 0
transform 1 0 10856 0 1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1546_
timestamp 0
transform 1 0 5152 0 1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1547_
timestamp 0
transform 1 0 9200 0 -1 23392
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1548_
timestamp 0
transform 1 0 11086 0 1 22848
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1549_
timestamp 0
transform 1 0 5520 0 1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1550_
timestamp 0
transform 1 0 8648 0 1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1551_
timestamp 0
transform 1 0 13800 0 1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1552_
timestamp 0
transform 1 0 14168 0 1 13600
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1553_
timestamp 0
transform 1 0 6348 0 -1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1554_
timestamp 0
transform 1 0 5888 0 1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1555_
timestamp 0
transform 1 0 7222 0 -1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1556_
timestamp 0
transform 1 0 12926 0 1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1557_
timestamp 0
transform 1 0 10810 0 1 10880
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1558_
timestamp 0
transform 1 0 5888 0 1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1559_
timestamp 0
transform 1 0 8648 0 1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1560_
timestamp 0
transform 1 0 10948 0 1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1561_
timestamp 0
transform 1 0 6670 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1562_
timestamp 0
transform 1 0 8510 0 1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1563_
timestamp 0
transform 1 0 12788 0 -1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1564_
timestamp 0
transform 1 0 12926 0 1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1565_
timestamp 0
transform 1 0 7268 0 -1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1566_
timestamp 0
transform 1 0 7222 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1567_
timestamp 0
transform 1 0 7406 0 1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1568_
timestamp 0
transform 1 0 12788 0 -1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1569_
timestamp 0
transform 1 0 10028 0 -1 15232
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1570_
timestamp 0
transform 1 0 7636 0 1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1571_
timestamp 0
transform 1 0 8234 0 1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1572_
timestamp 0
transform 1 0 11546 0 -1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1573_
timestamp 0
transform 1 0 7406 0 1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1574_
timestamp 0
transform 1 0 8648 0 1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1575_
timestamp 0
transform 1 0 13248 0 1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1576_
timestamp 0
transform 1 0 11408 0 1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1577_
timestamp 0
transform 1 0 3496 0 -1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1578_
timestamp 0
transform 1 0 3220 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1579_
timestamp 0
transform 1 0 4646 0 1 25568
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1580_
timestamp 0
transform 1 0 15180 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1581_
timestamp 0
transform 1 0 10580 0 1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1582_
timestamp 0
transform 1 0 5152 0 1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1583_
timestamp 0
transform 1 0 8188 0 1 24480
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1584_
timestamp 0
transform 1 0 9108 0 -1 22304
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1585_
timestamp 0
transform 1 0 3542 0 -1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1586_
timestamp 0
transform 1 0 8648 0 1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1587_
timestamp 0
transform 1 0 12926 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1588_
timestamp 0
transform 1 0 15548 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1589_
timestamp 0
transform 1 0 6164 0 -1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1590_
timestamp 0
transform 1 0 6578 0 -1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1591_
timestamp 0
transform 1 0 5520 0 1 24480
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1592_
timestamp 0
transform 1 0 15962 0 1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1593_
timestamp 0
transform 1 0 10948 0 1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1594_
timestamp 0
transform 1 0 5750 0 1 14144
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1595_
timestamp 0
transform 1 0 8786 0 -1 20128
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1596_
timestamp 0
transform 1 0 11638 0 -1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1597_
timestamp 0
transform 1 0 6670 0 -1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1598_
timestamp 0
transform 1 0 8648 0 1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1599_
timestamp 0
transform 1 0 15180 0 -1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1600_
timestamp 0
transform 1 0 12788 0 -1 11968
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1601_
timestamp 0
transform 1 0 3404 0 -1 22848
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1602_
timestamp 0
transform 1 0 3450 0 -1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1603_
timestamp 0
transform 1 0 3450 0 -1 23936
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1604_
timestamp 0
transform 1 0 16192 0 1 17952
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1605_
timestamp 0
transform 1 0 10764 0 1 15776
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1606_
timestamp 0
transform 1 0 4508 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1607_
timestamp 0
transform 1 0 8280 0 1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1608_
timestamp 0
transform 1 0 9660 0 -1 21760
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1609_
timestamp 0
transform 1 0 3404 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1610_
timestamp 0
transform 1 0 9108 0 -1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1611_
timestamp 0
transform 1 0 12696 0 -1 16320
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1612_
timestamp 0
transform 1 0 15778 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1613_
timestamp 0
transform 1 0 7268 0 -1 21216
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1614_
timestamp 0
transform 1 0 7222 0 -1 17408
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1615_
timestamp 0
transform 1 0 6900 0 -1 24480
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1616_
timestamp 0
transform 1 0 12972 0 1 19584
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1617_
timestamp 0
transform 1 0 10028 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1618_
timestamp 0
transform 1 0 6670 0 -1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1619_
timestamp 0
transform 1 0 8050 0 1 23936
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1620_
timestamp 0
transform 1 0 10810 0 1 20672
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1621_
timestamp 0
transform 1 0 7268 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1622_
timestamp 0
transform 1 0 8648 0 1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1623_
timestamp 0
transform 1 0 12788 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1624_
timestamp 0
transform 1 0 12374 0 -1 14688
box 0 -24 1104 296
use sky130_fd_sc_hd__dfrtp_1  _1625_
timestamp 0
transform 1 0 4784 0 1 28832
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_1  _1626_
timestamp 0
transform 1 0 4692 0 1 11968
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_1  _1627_
timestamp 0
transform 1 0 4692 0 -1 28832
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_1  _1628_
timestamp 0
transform 1 0 20194 0 -1 28288
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_4  _1629_
timestamp 0
transform 1 0 13524 0 1 10336
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1630_
timestamp 0
transform 1 0 4968 0 1 10336
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_4  _1631_
timestamp 0
transform 1 0 20286 0 -1 27200
box 0 -24 1058 296
use sky130_fd_sc_hd__dfrtp_1  _1632_
timestamp 0
transform 1 0 20148 0 -1 28832
box 0 -24 920 296
use sky130_fd_sc_hd__dfrtp_1  _1633_
timestamp 0
transform 1 0 5152 0 1 17952
box 0 -24 920 296
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 0
transform 1 0 18676 0 1 27744
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 0
transform 1 0 17204 0 1 28288
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 0
transform 1 0 11730 0 -1 26656
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 0
transform 1 0 13156 0 -1 29376
box 0 -24 736 296
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 0
transform 1 0 11270 0 1 26656
box 0 -24 736 296
use sky130_fd_sc_hd__edfxtp_1  _1639_
timestamp 0
transform 1 0 28290 0 -1 5984
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1640_
timestamp 0
transform 1 0 28382 0 -1 16864
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1641_
timestamp 0
transform 1 0 28198 0 -1 13056
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1642_
timestamp 0
transform 1 0 23276 0 -1 7616
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1643_
timestamp 0
transform 1 0 28382 0 -1 18496
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1644_
timestamp 0
transform 1 0 24380 0 1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1645_
timestamp 0
transform 1 0 17664 0 -1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1646_
timestamp 0
transform 1 0 21436 0 1 19040
box 0 -24 1104 296
use sky130_fd_sc_hd__edfxtp_1  _1647_
timestamp 0
transform 1 0 20470 0 -1 11424
box 0 -24 1104 296
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 0
transform 1 0 18676 0 -1 28288
box 0 -24 736 296
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform 1 0 8740 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 0
transform 1 0 14582 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__clkbuf_4  clkbuf_0_SysClk
timestamp 0
transform 1 0 8740 0 1 8160
box 0 -24 276 296
use sky130_fd_sc_hd__clkbuf_4  clkbuf_1_0__f_SysClk
timestamp 0
transform 1 0 7084 0 -1 7616
box 0 -24 276 296
use sky130_fd_sc_hd__clkbuf_4  clkbuf_1_1__f_SysClk
timestamp 0
transform 1 0 9430 0 -1 8704
box 0 -24 276 296
use sky130_fd_sc_hd__clkinv_2  clkload0
timestamp 0
transform 1 0 9292 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_0_0
timestamp 0
transform 1 0 3036 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_8
timestamp 0
transform 1 0 3404 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_16
timestamp 0
transform 1 0 3772 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_24
timestamp 0
transform 1 0 4140 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_0_28
timestamp 0
transform 1 0 4324 0 1 3264
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_0_31
timestamp 0
transform 1 0 4462 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_39
timestamp 0
transform 1 0 4830 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_47
timestamp 0
transform 1 0 5198 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_55
timestamp 0
transform 1 0 5566 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_59
timestamp 0
transform 1 0 5750 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_61
timestamp 0
transform 1 0 5842 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_69
timestamp 0
transform 1 0 6210 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_77
timestamp 0
transform 1 0 6578 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_85
timestamp 0
transform 1 0 6946 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 0
transform 1 0 7130 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_91
timestamp 0
transform 1 0 7222 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_99
timestamp 0
transform 1 0 7590 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_107
timestamp 0
transform 1 0 7958 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_115
timestamp 0
transform 1 0 8326 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 0
transform 1 0 8510 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_121
timestamp 0
transform 1 0 8602 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_129
timestamp 0
transform 1 0 8970 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_137
timestamp 0
transform 1 0 9338 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_145
timestamp 0
transform 1 0 9706 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 0
transform 1 0 9890 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_151
timestamp 0
transform 1 0 9982 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_159
timestamp 0
transform 1 0 10350 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_167
timestamp 0
transform 1 0 10718 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_175
timestamp 0
transform 1 0 11086 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_179
timestamp 0
transform 1 0 11270 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_181
timestamp 0
transform 1 0 11362 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_189
timestamp 0
transform 1 0 11730 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_197
timestamp 0
transform 1 0 12098 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_205
timestamp 0
transform 1 0 12466 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_209
timestamp 0
transform 1 0 12650 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_211
timestamp 0
transform 1 0 12742 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_219
timestamp 0
transform 1 0 13110 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_227
timestamp 0
transform 1 0 13478 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_235
timestamp 0
transform 1 0 13846 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_239
timestamp 0
transform 1 0 14030 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_241
timestamp 0
transform 1 0 14122 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_249
timestamp 0
transform 1 0 14490 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_257
timestamp 0
transform 1 0 14858 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_265
timestamp 0
transform 1 0 15226 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_269
timestamp 0
transform 1 0 15410 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_271
timestamp 0
transform 1 0 15502 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_279
timestamp 0
transform 1 0 15870 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_287
timestamp 0
transform 1 0 16238 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_295
timestamp 0
transform 1 0 16606 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_299
timestamp 0
transform 1 0 16790 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_301
timestamp 0
transform 1 0 16882 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_309
timestamp 0
transform 1 0 17250 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_317
timestamp 0
transform 1 0 17618 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_325
timestamp 0
transform 1 0 17986 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_329
timestamp 0
transform 1 0 18170 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_331
timestamp 0
transform 1 0 18262 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_339
timestamp 0
transform 1 0 18630 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_347
timestamp 0
transform 1 0 18998 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_355
timestamp 0
transform 1 0 19366 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_359
timestamp 0
transform 1 0 19550 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_361
timestamp 0
transform 1 0 19642 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_369
timestamp 0
transform 1 0 20010 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_377
timestamp 0
transform 1 0 20378 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_385
timestamp 0
transform 1 0 20746 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_389
timestamp 0
transform 1 0 20930 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_391
timestamp 0
transform 1 0 21022 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_399
timestamp 0
transform 1 0 21390 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_407
timestamp 0
transform 1 0 21758 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_415
timestamp 0
transform 1 0 22126 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 0
transform 1 0 22310 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_421
timestamp 0
transform 1 0 22402 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_429
timestamp 0
transform 1 0 22770 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_437
timestamp 0
transform 1 0 23138 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_445
timestamp 0
transform 1 0 23506 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_449
timestamp 0
transform 1 0 23690 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_451
timestamp 0
transform 1 0 23782 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_459
timestamp 0
transform 1 0 24150 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_467
timestamp 0
transform 1 0 24518 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_475
timestamp 0
transform 1 0 24886 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_479
timestamp 0
transform 1 0 25070 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_481
timestamp 0
transform 1 0 25162 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_489
timestamp 0
transform 1 0 25530 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_497
timestamp 0
transform 1 0 25898 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_505
timestamp 0
transform 1 0 26266 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_509
timestamp 0
transform 1 0 26450 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_511
timestamp 0
transform 1 0 26542 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_519
timestamp 0
transform 1 0 26910 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_527
timestamp 0
transform 1 0 27278 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_535
timestamp 0
transform 1 0 27646 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_539
timestamp 0
transform 1 0 27830 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_541
timestamp 0
transform 1 0 27922 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_549
timestamp 0
transform 1 0 28290 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_0_557
timestamp 0
transform 1 0 28658 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_565
timestamp 0
transform 1 0 29026 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_0_569
timestamp 0
transform 1 0 29210 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_0_571
timestamp 0
transform 1 0 29302 0 1 3264
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_0_579
timestamp 0
transform 1 0 29670 0 1 3264
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_0_583
timestamp 0
transform 1 0 29854 0 1 3264
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_0_585
timestamp 0
transform 1 0 29946 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_0
timestamp 0
transform 1 0 3036 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_8
timestamp 0
transform 1 0 3404 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_16
timestamp 0
transform 1 0 3772 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_24
timestamp 0
transform 1 0 4140 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_32
timestamp 0
transform 1 0 4508 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_40
timestamp 0
transform 1 0 4876 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_48
timestamp 0
transform 1 0 5244 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_1_56
timestamp 0
transform 1 0 5612 0 -1 3808
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_1_61
timestamp 0
transform 1 0 5842 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_69
timestamp 0
transform 1 0 6210 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_77
timestamp 0
transform 1 0 6578 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_85
timestamp 0
transform 1 0 6946 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_93
timestamp 0
transform 1 0 7314 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_101
timestamp 0
transform 1 0 7682 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_109
timestamp 0
transform 1 0 8050 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_117
timestamp 0
transform 1 0 8418 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 0
transform 1 0 8510 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_121
timestamp 0
transform 1 0 8602 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_129
timestamp 0
transform 1 0 8970 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_137
timestamp 0
transform 1 0 9338 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_145
timestamp 0
transform 1 0 9706 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_153
timestamp 0
transform 1 0 10074 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_161
timestamp 0
transform 1 0 10442 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_169
timestamp 0
transform 1 0 10810 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 0
transform 1 0 11178 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_179
timestamp 0
transform 1 0 11270 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_181
timestamp 0
transform 1 0 11362 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_189
timestamp 0
transform 1 0 11730 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_197
timestamp 0
transform 1 0 12098 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_205
timestamp 0
transform 1 0 12466 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_213
timestamp 0
transform 1 0 12834 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_221
timestamp 0
transform 1 0 13202 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_229
timestamp 0
transform 1 0 13570 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_237
timestamp 0
transform 1 0 13938 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_239
timestamp 0
transform 1 0 14030 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_241
timestamp 0
transform 1 0 14122 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_249
timestamp 0
transform 1 0 14490 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_257
timestamp 0
transform 1 0 14858 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_265
timestamp 0
transform 1 0 15226 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_273
timestamp 0
transform 1 0 15594 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_281
timestamp 0
transform 1 0 15962 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_289
timestamp 0
transform 1 0 16330 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 0
transform 1 0 16698 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_299
timestamp 0
transform 1 0 16790 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_301
timestamp 0
transform 1 0 16882 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_309
timestamp 0
transform 1 0 17250 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_317
timestamp 0
transform 1 0 17618 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_325
timestamp 0
transform 1 0 17986 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_333
timestamp 0
transform 1 0 18354 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_341
timestamp 0
transform 1 0 18722 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_349
timestamp 0
transform 1 0 19090 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_357
timestamp 0
transform 1 0 19458 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_359
timestamp 0
transform 1 0 19550 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_361
timestamp 0
transform 1 0 19642 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_369
timestamp 0
transform 1 0 20010 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_377
timestamp 0
transform 1 0 20378 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_385
timestamp 0
transform 1 0 20746 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_393
timestamp 0
transform 1 0 21114 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_401
timestamp 0
transform 1 0 21482 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_409
timestamp 0
transform 1 0 21850 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_417
timestamp 0
transform 1 0 22218 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_419
timestamp 0
transform 1 0 22310 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_421
timestamp 0
transform 1 0 22402 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_429
timestamp 0
transform 1 0 22770 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_437
timestamp 0
transform 1 0 23138 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_445
timestamp 0
transform 1 0 23506 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_453
timestamp 0
transform 1 0 23874 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_461
timestamp 0
transform 1 0 24242 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_469
timestamp 0
transform 1 0 24610 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_477
timestamp 0
transform 1 0 24978 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_479
timestamp 0
transform 1 0 25070 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_481
timestamp 0
transform 1 0 25162 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_489
timestamp 0
transform 1 0 25530 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_497
timestamp 0
transform 1 0 25898 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_505
timestamp 0
transform 1 0 26266 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_513
timestamp 0
transform 1 0 26634 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_521
timestamp 0
transform 1 0 27002 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_529
timestamp 0
transform 1 0 27370 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_1_537
timestamp 0
transform 1 0 27738 0 -1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_1_539
timestamp 0
transform 1 0 27830 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_1_541
timestamp 0
transform 1 0 27922 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_549
timestamp 0
transform 1 0 28290 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_557
timestamp 0
transform 1 0 28658 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_565
timestamp 0
transform 1 0 29026 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_1_573
timestamp 0
transform 1 0 29394 0 -1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_1_581
timestamp 0
transform 1 0 29762 0 -1 3808
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_1_585
timestamp 0
transform 1 0 29946 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_0
timestamp 0
transform 1 0 3036 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_8
timestamp 0
transform 1 0 3404 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_16
timestamp 0
transform 1 0 3772 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_2_24
timestamp 0
transform 1 0 4140 0 1 3808
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_2_28
timestamp 0
transform 1 0 4324 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_2_31
timestamp 0
transform 1 0 4462 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_39
timestamp 0
transform 1 0 4830 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_47
timestamp 0
transform 1 0 5198 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_55
timestamp 0
transform 1 0 5566 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_63
timestamp 0
transform 1 0 5934 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_71
timestamp 0
transform 1 0 6302 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_79
timestamp 0
transform 1 0 6670 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_87
timestamp 0
transform 1 0 7038 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 0
transform 1 0 7130 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_91
timestamp 0
transform 1 0 7222 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_99
timestamp 0
transform 1 0 7590 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_107
timestamp 0
transform 1 0 7958 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_115
timestamp 0
transform 1 0 8326 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_123
timestamp 0
transform 1 0 8694 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_131
timestamp 0
transform 1 0 9062 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_139
timestamp 0
transform 1 0 9430 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp 0
transform 1 0 9798 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 0
transform 1 0 9890 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_151
timestamp 0
transform 1 0 9982 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_159
timestamp 0
transform 1 0 10350 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_167
timestamp 0
transform 1 0 10718 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_175
timestamp 0
transform 1 0 11086 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_183
timestamp 0
transform 1 0 11454 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_191
timestamp 0
transform 1 0 11822 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_199
timestamp 0
transform 1 0 12190 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_207
timestamp 0
transform 1 0 12558 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_209
timestamp 0
transform 1 0 12650 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_211
timestamp 0
transform 1 0 12742 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_219
timestamp 0
transform 1 0 13110 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_227
timestamp 0
transform 1 0 13478 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_235
timestamp 0
transform 1 0 13846 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_243
timestamp 0
transform 1 0 14214 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_251
timestamp 0
transform 1 0 14582 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_259
timestamp 0
transform 1 0 14950 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_267
timestamp 0
transform 1 0 15318 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_269
timestamp 0
transform 1 0 15410 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_271
timestamp 0
transform 1 0 15502 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_279
timestamp 0
transform 1 0 15870 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_287
timestamp 0
transform 1 0 16238 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_295
timestamp 0
transform 1 0 16606 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_303
timestamp 0
transform 1 0 16974 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_311
timestamp 0
transform 1 0 17342 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_319
timestamp 0
transform 1 0 17710 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_327
timestamp 0
transform 1 0 18078 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_329
timestamp 0
transform 1 0 18170 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_2_331
timestamp 0
transform 1 0 18262 0 1 3808
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_2_335
timestamp 0
transform 1 0 18446 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_2_350
timestamp 0
transform 1 0 19136 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_358
timestamp 0
transform 1 0 19504 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_366
timestamp 0
transform 1 0 19872 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_374
timestamp 0
transform 1 0 20240 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_382
timestamp 0
transform 1 0 20608 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_391
timestamp 0
transform 1 0 21022 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_399
timestamp 0
transform 1 0 21390 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_407
timestamp 0
transform 1 0 21758 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_415
timestamp 0
transform 1 0 22126 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_423
timestamp 0
transform 1 0 22494 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_431
timestamp 0
transform 1 0 22862 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_439
timestamp 0
transform 1 0 23230 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_447
timestamp 0
transform 1 0 23598 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_449
timestamp 0
transform 1 0 23690 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_451
timestamp 0
transform 1 0 23782 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_459
timestamp 0
transform 1 0 24150 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_467
timestamp 0
transform 1 0 24518 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_475
timestamp 0
transform 1 0 24886 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_483
timestamp 0
transform 1 0 25254 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_491
timestamp 0
transform 1 0 25622 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_499
timestamp 0
transform 1 0 25990 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_507
timestamp 0
transform 1 0 26358 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_509
timestamp 0
transform 1 0 26450 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_511
timestamp 0
transform 1 0 26542 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_519
timestamp 0
transform 1 0 26910 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_527
timestamp 0
transform 1 0 27278 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_535
timestamp 0
transform 1 0 27646 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_543
timestamp 0
transform 1 0 28014 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_551
timestamp 0
transform 1 0 28382 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_2_559
timestamp 0
transform 1 0 28750 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_2_567
timestamp 0
transform 1 0 29118 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_569
timestamp 0
transform 1 0 29210 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_2_571
timestamp 0
transform 1 0 29302 0 1 3808
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_2_579
timestamp 0
transform 1 0 29670 0 1 3808
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_2_583
timestamp 0
transform 1 0 29854 0 1 3808
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_2_585
timestamp 0
transform 1 0 29946 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_0
timestamp 0
transform 1 0 3036 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_8
timestamp 0
transform 1 0 3404 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_16
timestamp 0
transform 1 0 3772 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_24
timestamp 0
transform 1 0 4140 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_32
timestamp 0
transform 1 0 4508 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_40
timestamp 0
transform 1 0 4876 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_48
timestamp 0
transform 1 0 5244 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_3_56
timestamp 0
transform 1 0 5612 0 -1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_3_61
timestamp 0
transform 1 0 5842 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_69
timestamp 0
transform 1 0 6210 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_77
timestamp 0
transform 1 0 6578 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_85
timestamp 0
transform 1 0 6946 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_93
timestamp 0
transform 1 0 7314 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_101
timestamp 0
transform 1 0 7682 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_109
timestamp 0
transform 1 0 8050 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 0
transform 1 0 8418 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 0
transform 1 0 8510 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_121
timestamp 0
transform 1 0 8602 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_129
timestamp 0
transform 1 0 8970 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_137
timestamp 0
transform 1 0 9338 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_145
timestamp 0
transform 1 0 9706 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_153
timestamp 0
transform 1 0 10074 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_161
timestamp 0
transform 1 0 10442 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_169
timestamp 0
transform 1 0 10810 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_177
timestamp 0
transform 1 0 11178 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_179
timestamp 0
transform 1 0 11270 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_181
timestamp 0
transform 1 0 11362 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_189
timestamp 0
transform 1 0 11730 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_197
timestamp 0
transform 1 0 12098 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_205
timestamp 0
transform 1 0 12466 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_213
timestamp 0
transform 1 0 12834 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_221
timestamp 0
transform 1 0 13202 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_229
timestamp 0
transform 1 0 13570 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_237
timestamp 0
transform 1 0 13938 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_239
timestamp 0
transform 1 0 14030 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_241
timestamp 0
transform 1 0 14122 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_249
timestamp 0
transform 1 0 14490 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_257
timestamp 0
transform 1 0 14858 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_265
timestamp 0
transform 1 0 15226 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_273
timestamp 0
transform 1 0 15594 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_281
timestamp 0
transform 1 0 15962 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_289
timestamp 0
transform 1 0 16330 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 0
transform 1 0 16698 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_299
timestamp 0
transform 1 0 16790 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_301
timestamp 0
transform 1 0 16882 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_309
timestamp 0
transform 1 0 17250 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_317
timestamp 0
transform 1 0 17618 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_325
timestamp 0
transform 1 0 17986 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_333
timestamp 0
transform 1 0 18354 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_341
timestamp 0
transform 1 0 18722 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_349
timestamp 0
transform 1 0 19090 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_357
timestamp 0
transform 1 0 19458 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_359
timestamp 0
transform 1 0 19550 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_361
timestamp 0
transform 1 0 19642 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_369
timestamp 0
transform 1 0 20010 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_377
timestamp 0
transform 1 0 20378 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_385
timestamp 0
transform 1 0 20746 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_393
timestamp 0
transform 1 0 21114 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_401
timestamp 0
transform 1 0 21482 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_409
timestamp 0
transform 1 0 21850 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_417
timestamp 0
transform 1 0 22218 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_419
timestamp 0
transform 1 0 22310 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_421
timestamp 0
transform 1 0 22402 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_429
timestamp 0
transform 1 0 22770 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_437
timestamp 0
transform 1 0 23138 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_445
timestamp 0
transform 1 0 23506 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_453
timestamp 0
transform 1 0 23874 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_461
timestamp 0
transform 1 0 24242 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_469
timestamp 0
transform 1 0 24610 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_477
timestamp 0
transform 1 0 24978 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_479
timestamp 0
transform 1 0 25070 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_481
timestamp 0
transform 1 0 25162 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_489
timestamp 0
transform 1 0 25530 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_497
timestamp 0
transform 1 0 25898 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_505
timestamp 0
transform 1 0 26266 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_513
timestamp 0
transform 1 0 26634 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_521
timestamp 0
transform 1 0 27002 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_529
timestamp 0
transform 1 0 27370 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_3_537
timestamp 0
transform 1 0 27738 0 -1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_3_539
timestamp 0
transform 1 0 27830 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_3_541
timestamp 0
transform 1 0 27922 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_549
timestamp 0
transform 1 0 28290 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_557
timestamp 0
transform 1 0 28658 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_565
timestamp 0
transform 1 0 29026 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_3_573
timestamp 0
transform 1 0 29394 0 -1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_3_581
timestamp 0
transform 1 0 29762 0 -1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_3_585
timestamp 0
transform 1 0 29946 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_0
timestamp 0
transform 1 0 3036 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_8
timestamp 0
transform 1 0 3404 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_16
timestamp 0
transform 1 0 3772 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_4_24
timestamp 0
transform 1 0 4140 0 1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_4_28
timestamp 0
transform 1 0 4324 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_4_31
timestamp 0
transform 1 0 4462 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_39
timestamp 0
transform 1 0 4830 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_47
timestamp 0
transform 1 0 5198 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_55
timestamp 0
transform 1 0 5566 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_63
timestamp 0
transform 1 0 5934 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_71
timestamp 0
transform 1 0 6302 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_79
timestamp 0
transform 1 0 6670 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 0
transform 1 0 7038 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 0
transform 1 0 7130 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_91
timestamp 0
transform 1 0 7222 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_99
timestamp 0
transform 1 0 7590 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_107
timestamp 0
transform 1 0 7958 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_115
timestamp 0
transform 1 0 8326 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_123
timestamp 0
transform 1 0 8694 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_131
timestamp 0
transform 1 0 9062 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_139
timestamp 0
transform 1 0 9430 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_4_147
timestamp 0
transform 1 0 9798 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_149
timestamp 0
transform 1 0 9890 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_151
timestamp 0
transform 1 0 9982 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_159
timestamp 0
transform 1 0 10350 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_167
timestamp 0
transform 1 0 10718 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_175
timestamp 0
transform 1 0 11086 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_183
timestamp 0
transform 1 0 11454 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_191
timestamp 0
transform 1 0 11822 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_199
timestamp 0
transform 1 0 12190 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_4_207
timestamp 0
transform 1 0 12558 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 0
transform 1 0 12650 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_211
timestamp 0
transform 1 0 12742 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_219
timestamp 0
transform 1 0 13110 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_227
timestamp 0
transform 1 0 13478 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_235
timestamp 0
transform 1 0 13846 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_243
timestamp 0
transform 1 0 14214 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_251
timestamp 0
transform 1 0 14582 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_259
timestamp 0
transform 1 0 14950 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_4_267
timestamp 0
transform 1 0 15318 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_269
timestamp 0
transform 1 0 15410 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_271
timestamp 0
transform 1 0 15502 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_279
timestamp 0
transform 1 0 15870 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_4_287
timestamp 0
transform 1 0 16238 0 1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_4_291
timestamp 0
transform 1 0 16422 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_293
timestamp 0
transform 1 0 16514 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_310
timestamp 0
transform 1 0 17296 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_318
timestamp 0
transform 1 0 17664 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_4_326
timestamp 0
transform 1 0 18032 0 1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_4_331
timestamp 0
transform 1 0 18262 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_339
timestamp 0
transform 1 0 18630 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_347
timestamp 0
transform 1 0 18998 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_355
timestamp 0
transform 1 0 19366 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_363
timestamp 0
transform 1 0 19734 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_371
timestamp 0
transform 1 0 20102 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_379
timestamp 0
transform 1 0 20470 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_4_387
timestamp 0
transform 1 0 20838 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_389
timestamp 0
transform 1 0 20930 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_391
timestamp 0
transform 1 0 21022 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_399
timestamp 0
transform 1 0 21390 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_407
timestamp 0
transform 1 0 21758 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_415
timestamp 0
transform 1 0 22126 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_423
timestamp 0
transform 1 0 22494 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_431
timestamp 0
transform 1 0 22862 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_439
timestamp 0
transform 1 0 23230 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_4_447
timestamp 0
transform 1 0 23598 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_449
timestamp 0
transform 1 0 23690 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_4_451
timestamp 0
transform 1 0 23782 0 1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_4_455
timestamp 0
transform 1 0 23966 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_4_481
timestamp 0
transform 1 0 25162 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_489
timestamp 0
transform 1 0 25530 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_497
timestamp 0
transform 1 0 25898 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_4_505
timestamp 0
transform 1 0 26266 0 1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_4_509
timestamp 0
transform 1 0 26450 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_511
timestamp 0
transform 1 0 26542 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_519
timestamp 0
transform 1 0 26910 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_527
timestamp 0
transform 1 0 27278 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_535
timestamp 0
transform 1 0 27646 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_543
timestamp 0
transform 1 0 28014 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_551
timestamp 0
transform 1 0 28382 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_4_559
timestamp 0
transform 1 0 28750 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_4_567
timestamp 0
transform 1 0 29118 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_569
timestamp 0
transform 1 0 29210 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_4_571
timestamp 0
transform 1 0 29302 0 1 4352
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_4_579
timestamp 0
transform 1 0 29670 0 1 4352
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_4_583
timestamp 0
transform 1 0 29854 0 1 4352
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_4_585
timestamp 0
transform 1 0 29946 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_5_0
timestamp 0
transform 1 0 3036 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_8
timestamp 0
transform 1 0 3404 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_16
timestamp 0
transform 1 0 3772 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_24
timestamp 0
transform 1 0 4140 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_32
timestamp 0
transform 1 0 4508 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_40
timestamp 0
transform 1 0 4876 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_48
timestamp 0
transform 1 0 5244 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_5_56
timestamp 0
transform 1 0 5612 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_5_61
timestamp 0
transform 1 0 5842 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_69
timestamp 0
transform 1 0 6210 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_77
timestamp 0
transform 1 0 6578 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_85
timestamp 0
transform 1 0 6946 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_93
timestamp 0
transform 1 0 7314 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_101
timestamp 0
transform 1 0 7682 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_109
timestamp 0
transform 1 0 8050 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_5_117
timestamp 0
transform 1 0 8418 0 -1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp 0
transform 1 0 8510 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_5_121
timestamp 0
transform 1 0 8602 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_129
timestamp 0
transform 1 0 8970 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_137
timestamp 0
transform 1 0 9338 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_145
timestamp 0
transform 1 0 9706 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_153
timestamp 0
transform 1 0 10074 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_161
timestamp 0
transform 1 0 10442 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_169
timestamp 0
transform 1 0 10810 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 0
transform 1 0 11178 0 -1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_5_179
timestamp 0
transform 1 0 11270 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_5_181
timestamp 0
transform 1 0 11362 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_189
timestamp 0
transform 1 0 11730 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_197
timestamp 0
transform 1 0 12098 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_205
timestamp 0
transform 1 0 12466 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_213
timestamp 0
transform 1 0 12834 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_221
timestamp 0
transform 1 0 13202 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_229
timestamp 0
transform 1 0 13570 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_5_237
timestamp 0
transform 1 0 13938 0 -1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_5_239
timestamp 0
transform 1 0 14030 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_5_241
timestamp 0
transform 1 0 14122 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_249
timestamp 0
transform 1 0 14490 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_257
timestamp 0
transform 1 0 14858 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_265
timestamp 0
transform 1 0 15226 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_273
timestamp 0
transform 1 0 15594 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_281
timestamp 0
transform 1 0 15962 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_5_289
timestamp 0
transform 1 0 16330 0 -1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_5_295
timestamp 0
transform 1 0 16606 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_5_299
timestamp 0
transform 1 0 16790 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_5_301
timestamp 0
transform 1 0 16882 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_5_309
timestamp 0
transform 1 0 17250 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_317
timestamp 0
transform 1 0 17618 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_325
timestamp 0
transform 1 0 17986 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_5_333
timestamp 0
transform 1 0 18354 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_5_350
timestamp 0
transform 1 0 19136 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_5_358
timestamp 0
transform 1 0 19504 0 -1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_5_361
timestamp 0
transform 1 0 19642 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_5_376
timestamp 0
transform 1 0 20332 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_384
timestamp 0
transform 1 0 20700 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_5_416
timestamp 0
transform 1 0 22172 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_5_421
timestamp 0
transform 1 0 22402 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_429
timestamp 0
transform 1 0 22770 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_437
timestamp 0
transform 1 0 23138 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_445
timestamp 0
transform 1 0 23506 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_453
timestamp 0
transform 1 0 23874 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_461
timestamp 0
transform 1 0 24242 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_469
timestamp 0
transform 1 0 24610 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_5_477
timestamp 0
transform 1 0 24978 0 -1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_5_479
timestamp 0
transform 1 0 25070 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_5_481
timestamp 0
transform 1 0 25162 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_489
timestamp 0
transform 1 0 25530 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_497
timestamp 0
transform 1 0 25898 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_505
timestamp 0
transform 1 0 26266 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_513
timestamp 0
transform 1 0 26634 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_521
timestamp 0
transform 1 0 27002 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_529
timestamp 0
transform 1 0 27370 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_5_537
timestamp 0
transform 1 0 27738 0 -1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_5_539
timestamp 0
transform 1 0 27830 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_5_541
timestamp 0
transform 1 0 27922 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_549
timestamp 0
transform 1 0 28290 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_557
timestamp 0
transform 1 0 28658 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_565
timestamp 0
transform 1 0 29026 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_5_573
timestamp 0
transform 1 0 29394 0 -1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_5_581
timestamp 0
transform 1 0 29762 0 -1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_5_585
timestamp 0
transform 1 0 29946 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_0
timestamp 0
transform 1 0 3036 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_8
timestamp 0
transform 1 0 3404 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_16
timestamp 0
transform 1 0 3772 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_6_24
timestamp 0
transform 1 0 4140 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_6_28
timestamp 0
transform 1 0 4324 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_6_31
timestamp 0
transform 1 0 4462 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_39
timestamp 0
transform 1 0 4830 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_47
timestamp 0
transform 1 0 5198 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_55
timestamp 0
transform 1 0 5566 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_63
timestamp 0
transform 1 0 5934 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_71
timestamp 0
transform 1 0 6302 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_79
timestamp 0
transform 1 0 6670 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 0
transform 1 0 7038 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 0
transform 1 0 7130 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_91
timestamp 0
transform 1 0 7222 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_99
timestamp 0
transform 1 0 7590 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_6_107
timestamp 0
transform 1 0 7958 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_109
timestamp 0
transform 1 0 8050 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_113
timestamp 0
transform 1 0 8234 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_121
timestamp 0
transform 1 0 8602 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_129
timestamp 0
transform 1 0 8970 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_137
timestamp 0
transform 1 0 9338 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_6_145
timestamp 0
transform 1 0 9706 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_6_149
timestamp 0
transform 1 0 9890 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_151
timestamp 0
transform 1 0 9982 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_159
timestamp 0
transform 1 0 10350 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_167
timestamp 0
transform 1 0 10718 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_175
timestamp 0
transform 1 0 11086 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_183
timestamp 0
transform 1 0 11454 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_191
timestamp 0
transform 1 0 11822 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_199
timestamp 0
transform 1 0 12190 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_6_207
timestamp 0
transform 1 0 12558 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_209
timestamp 0
transform 1 0 12650 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_211
timestamp 0
transform 1 0 12742 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_219
timestamp 0
transform 1 0 13110 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_227
timestamp 0
transform 1 0 13478 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_235
timestamp 0
transform 1 0 13846 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_243
timestamp 0
transform 1 0 14214 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_251
timestamp 0
transform 1 0 14582 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_259
timestamp 0
transform 1 0 14950 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_6_267
timestamp 0
transform 1 0 15318 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_269
timestamp 0
transform 1 0 15410 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_271
timestamp 0
transform 1 0 15502 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_279
timestamp 0
transform 1 0 15870 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_287
timestamp 0
transform 1 0 16238 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_295
timestamp 0
transform 1 0 16606 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_303
timestamp 0
transform 1 0 16974 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_311
timestamp 0
transform 1 0 17342 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_319
timestamp 0
transform 1 0 17710 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_6_327
timestamp 0
transform 1 0 18078 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_329
timestamp 0
transform 1 0 18170 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_6_331
timestamp 0
transform 1 0 18262 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_6_340
timestamp 0
transform 1 0 18676 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_348
timestamp 0
transform 1 0 19044 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_6_356
timestamp 0
transform 1 0 19412 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_6_371
timestamp 0
transform 1 0 20102 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_379
timestamp 0
transform 1 0 20470 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_6_387
timestamp 0
transform 1 0 20838 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_389
timestamp 0
transform 1 0 20930 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_6_391
timestamp 0
transform 1 0 21022 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_6_419
timestamp 0
transform 1 0 22310 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_427
timestamp 0
transform 1 0 22678 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_435
timestamp 0
transform 1 0 23046 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_6_443
timestamp 0
transform 1 0 23414 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_6_447
timestamp 0
transform 1 0 23598 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_449
timestamp 0
transform 1 0 23690 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_6_451
timestamp 0
transform 1 0 23782 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_6_479
timestamp 0
transform 1 0 25070 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_487
timestamp 0
transform 1 0 25438 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_495
timestamp 0
transform 1 0 25806 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_6_503
timestamp 0
transform 1 0 26174 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_6_507
timestamp 0
transform 1 0 26358 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_509
timestamp 0
transform 1 0 26450 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_511
timestamp 0
transform 1 0 26542 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_519
timestamp 0
transform 1 0 26910 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_527
timestamp 0
transform 1 0 27278 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_535
timestamp 0
transform 1 0 27646 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_543
timestamp 0
transform 1 0 28014 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_551
timestamp 0
transform 1 0 28382 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_6_559
timestamp 0
transform 1 0 28750 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_6_567
timestamp 0
transform 1 0 29118 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_569
timestamp 0
transform 1 0 29210 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_6_571
timestamp 0
transform 1 0 29302 0 1 4896
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_6_579
timestamp 0
transform 1 0 29670 0 1 4896
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_6_583
timestamp 0
transform 1 0 29854 0 1 4896
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_6_585
timestamp 0
transform 1 0 29946 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_7_0
timestamp 0
transform 1 0 3036 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_8
timestamp 0
transform 1 0 3404 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_16
timestamp 0
transform 1 0 3772 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_24
timestamp 0
transform 1 0 4140 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_32
timestamp 0
transform 1 0 4508 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_40
timestamp 0
transform 1 0 4876 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_48
timestamp 0
transform 1 0 5244 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_7_56
timestamp 0
transform 1 0 5612 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_7_61
timestamp 0
transform 1 0 5842 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_69
timestamp 0
transform 1 0 6210 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_77
timestamp 0
transform 1 0 6578 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_85
timestamp 0
transform 1 0 6946 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_93
timestamp 0
transform 1 0 7314 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 0
transform 1 0 7682 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_7_108
timestamp 0
transform 1 0 8004 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_7_115
timestamp 0
transform 1 0 8326 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 0
transform 1 0 8510 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_7_121
timestamp 0
transform 1 0 8602 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp 0
transform 1 0 8786 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 0
transform 1 0 8878 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_7_133
timestamp 0
transform 1 0 9154 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_141
timestamp 0
transform 1 0 9522 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 0
transform 1 0 9890 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_7_151
timestamp 0
transform 1 0 9982 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_7_155
timestamp 0
transform 1 0 10166 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_163
timestamp 0
transform 1 0 10534 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_171
timestamp 0
transform 1 0 10902 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_7_179
timestamp 0
transform 1 0 11270 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_7_181
timestamp 0
transform 1 0 11362 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_189
timestamp 0
transform 1 0 11730 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_197
timestamp 0
transform 1 0 12098 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_205
timestamp 0
transform 1 0 12466 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_213
timestamp 0
transform 1 0 12834 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_221
timestamp 0
transform 1 0 13202 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_229
timestamp 0
transform 1 0 13570 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_7_237
timestamp 0
transform 1 0 13938 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_7_239
timestamp 0
transform 1 0 14030 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_7_241
timestamp 0
transform 1 0 14122 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_249
timestamp 0
transform 1 0 14490 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_7_257
timestamp 0
transform 1 0 14858 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_7_259
timestamp 0
transform 1 0 14950 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_7_276
timestamp 0
transform 1 0 15732 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_7_285
timestamp 0
transform 1 0 16146 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_7_293
timestamp 0
transform 1 0 16514 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 0
transform 1 0 16698 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_7_299
timestamp 0
transform 1 0 16790 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_7_301
timestamp 0
transform 1 0 16882 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_7_309
timestamp 0
transform 1 0 17250 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_7_314
timestamp 0
transform 1 0 17480 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_322
timestamp 0
transform 1 0 17848 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_7_330
timestamp 0
transform 1 0 18216 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_7_336
timestamp 0
transform 1 0 18492 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_344
timestamp 0
transform 1 0 18860 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_352
timestamp 0
transform 1 0 19228 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_7_361
timestamp 0
transform 1 0 19642 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_7_365
timestamp 0
transform 1 0 19826 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_7_376
timestamp 0
transform 1 0 20332 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_384
timestamp 0
transform 1 0 20700 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_7_416
timestamp 0
transform 1 0 22172 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_7_421
timestamp 0
transform 1 0 22402 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_429
timestamp 0
transform 1 0 22770 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_437
timestamp 0
transform 1 0 23138 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_7_445
timestamp 0
transform 1 0 23506 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp 0
transform 1 0 23690 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_7_475
timestamp 0
transform 1 0 24886 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_7_479
timestamp 0
transform 1 0 25070 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_7_481
timestamp 0
transform 1 0 25162 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_7_493
timestamp 0
transform 1 0 25714 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_501
timestamp 0
transform 1 0 26082 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_509
timestamp 0
transform 1 0 26450 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_517
timestamp 0
transform 1 0 26818 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_525
timestamp 0
transform 1 0 27186 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_7_533
timestamp 0
transform 1 0 27554 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_7_537
timestamp 0
transform 1 0 27738 0 -1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_7_539
timestamp 0
transform 1 0 27830 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_7_541
timestamp 0
transform 1 0 27922 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_549
timestamp 0
transform 1 0 28290 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_557
timestamp 0
transform 1 0 28658 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_565
timestamp 0
transform 1 0 29026 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_7_573
timestamp 0
transform 1 0 29394 0 -1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_7_581
timestamp 0
transform 1 0 29762 0 -1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_7_585
timestamp 0
transform 1 0 29946 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_0
timestamp 0
transform 1 0 3036 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_8
timestamp 0
transform 1 0 3404 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_16
timestamp 0
transform 1 0 3772 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_8_24
timestamp 0
transform 1 0 4140 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_8_28
timestamp 0
transform 1 0 4324 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_8_31
timestamp 0
transform 1 0 4462 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_39
timestamp 0
transform 1 0 4830 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_47
timestamp 0
transform 1 0 5198 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_55
timestamp 0
transform 1 0 5566 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_63
timestamp 0
transform 1 0 5934 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_71
timestamp 0
transform 1 0 6302 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_79
timestamp 0
transform 1 0 6670 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 0
transform 1 0 7038 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 0
transform 1 0 7130 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_91
timestamp 0
transform 1 0 7222 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_99
timestamp 0
transform 1 0 7590 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 0
transform 1 0 7682 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_109
timestamp 0
transform 1 0 8050 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 0
transform 1 0 8418 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_8_124
timestamp 0
transform 1 0 8740 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_8_132
timestamp 0
transform 1 0 9108 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_140
timestamp 0
transform 1 0 9476 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 0
transform 1 0 9844 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_8_151
timestamp 0
transform 1 0 9982 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_8_159
timestamp 0
transform 1 0 10350 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_167
timestamp 0
transform 1 0 10718 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_175
timestamp 0
transform 1 0 11086 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_183
timestamp 0
transform 1 0 11454 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_191
timestamp 0
transform 1 0 11822 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_199
timestamp 0
transform 1 0 12190 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_207
timestamp 0
transform 1 0 12558 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_209
timestamp 0
transform 1 0 12650 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_211
timestamp 0
transform 1 0 12742 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_219
timestamp 0
transform 1 0 13110 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_227
timestamp 0
transform 1 0 13478 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_235
timestamp 0
transform 1 0 13846 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_243
timestamp 0
transform 1 0 14214 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_251
timestamp 0
transform 1 0 14582 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_259
timestamp 0
transform 1 0 14950 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_267
timestamp 0
transform 1 0 15318 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_269
timestamp 0
transform 1 0 15410 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_8_271
timestamp 0
transform 1 0 15502 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_8_279
timestamp 0
transform 1 0 15870 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_287
timestamp 0
transform 1 0 16238 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_8_295
timestamp 0
transform 1 0 16606 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_8_299
timestamp 0
transform 1 0 16790 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_8_304
timestamp 0
transform 1 0 17020 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_8_308
timestamp 0
transform 1 0 17204 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_8_325
timestamp 0
transform 1 0 17986 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_8_329
timestamp 0
transform 1 0 18170 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_8_331
timestamp 0
transform 1 0 18262 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_8_341
timestamp 0
transform 1 0 18722 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_349
timestamp 0
transform 1 0 19090 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_8_357
timestamp 0
transform 1 0 19458 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_8_361
timestamp 0
transform 1 0 19642 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 0
transform 1 0 19734 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_373
timestamp 0
transform 1 0 20194 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_381
timestamp 0
transform 1 0 20562 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_8_389
timestamp 0
transform 1 0 20930 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_391
timestamp 0
transform 1 0 21022 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_399
timestamp 0
transform 1 0 21390 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_407
timestamp 0
transform 1 0 21758 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_423
timestamp 0
transform 1 0 22494 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_431
timestamp 0
transform 1 0 22862 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_439
timestamp 0
transform 1 0 23230 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_447
timestamp 0
transform 1 0 23598 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_449
timestamp 0
transform 1 0 23690 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_451
timestamp 0
transform 1 0 23782 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_459
timestamp 0
transform 1 0 24150 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_467
timestamp 0
transform 1 0 24518 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_475
timestamp 0
transform 1 0 24886 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_483
timestamp 0
transform 1 0 25254 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_491
timestamp 0
transform 1 0 25622 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_499
timestamp 0
transform 1 0 25990 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_507
timestamp 0
transform 1 0 26358 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_509
timestamp 0
transform 1 0 26450 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_8_511
timestamp 0
transform 1 0 26542 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_8_520
timestamp 0
transform 1 0 26956 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_8_524
timestamp 0
transform 1 0 27140 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_8_528
timestamp 0
transform 1 0 27324 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_536
timestamp 0
transform 1 0 27692 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_544
timestamp 0
transform 1 0 28060 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_552
timestamp 0
transform 1 0 28428 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_8_560
timestamp 0
transform 1 0 28796 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_8_568
timestamp 0
transform 1 0 29164 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_8_571
timestamp 0
transform 1 0 29302 0 1 5440
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_8_579
timestamp 0
transform 1 0 29670 0 1 5440
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_8_583
timestamp 0
transform 1 0 29854 0 1 5440
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_8_585
timestamp 0
transform 1 0 29946 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_9_0
timestamp 0
transform 1 0 3036 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_8
timestamp 0
transform 1 0 3404 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_16
timestamp 0
transform 1 0 3772 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_24
timestamp 0
transform 1 0 4140 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_32
timestamp 0
transform 1 0 4508 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_40
timestamp 0
transform 1 0 4876 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_48
timestamp 0
transform 1 0 5244 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_56
timestamp 0
transform 1 0 5612 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_9_61
timestamp 0
transform 1 0 5842 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_69
timestamp 0
transform 1 0 6210 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_77
timestamp 0
transform 1 0 6578 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_85
timestamp 0
transform 1 0 6946 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_93
timestamp 0
transform 1 0 7314 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_104
timestamp 0
transform 1 0 7820 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_9_108
timestamp 0
transform 1 0 8004 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_9_116
timestamp 0
transform 1 0 8372 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_9_121
timestamp 0
transform 1 0 8602 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_129
timestamp 0
transform 1 0 8970 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_9_133
timestamp 0
transform 1 0 9154 0 -1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_9_135
timestamp 0
transform 1 0 9246 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_9_144
timestamp 0
transform 1 0 9660 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_9_158
timestamp 0
transform 1 0 10304 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_166
timestamp 0
transform 1 0 10672 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 0
transform 1 0 10856 0 -1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_9_176
timestamp 0
transform 1 0 11132 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_9_181
timestamp 0
transform 1 0 11362 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_9_189
timestamp 0
transform 1 0 11730 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_197
timestamp 0
transform 1 0 12098 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_205
timestamp 0
transform 1 0 12466 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_213
timestamp 0
transform 1 0 12834 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_221
timestamp 0
transform 1 0 13202 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_229
timestamp 0
transform 1 0 13570 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_9_237
timestamp 0
transform 1 0 13938 0 -1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_9_239
timestamp 0
transform 1 0 14030 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_9_241
timestamp 0
transform 1 0 14122 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_249
timestamp 0
transform 1 0 14490 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_257
timestamp 0
transform 1 0 14858 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_265
timestamp 0
transform 1 0 15226 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_273
timestamp 0
transform 1 0 15594 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_281
timestamp 0
transform 1 0 15962 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_289
timestamp 0
transform 1 0 16330 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_9_297
timestamp 0
transform 1 0 16698 0 -1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_9_299
timestamp 0
transform 1 0 16790 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_9_301
timestamp 0
transform 1 0 16882 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_9_312
timestamp 0
transform 1 0 17388 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_320
timestamp 0
transform 1 0 17756 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_328
timestamp 0
transform 1 0 18124 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_9_332
timestamp 0
transform 1 0 18308 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_9_347
timestamp 0
transform 1 0 18998 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_355
timestamp 0
transform 1 0 19366 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_9_359
timestamp 0
transform 1 0 19550 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_9_361
timestamp 0
transform 1 0 19642 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_9_374
timestamp 0
transform 1 0 20240 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_382
timestamp 0
transform 1 0 20608 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_390
timestamp 0
transform 1 0 20976 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_398
timestamp 0
transform 1 0 21344 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_406
timestamp 0
transform 1 0 21712 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_414
timestamp 0
transform 1 0 22080 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_9_418
timestamp 0
transform 1 0 22264 0 -1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_9_421
timestamp 0
transform 1 0 22402 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_429
timestamp 0
transform 1 0 22770 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_437
timestamp 0
transform 1 0 23138 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_445
timestamp 0
transform 1 0 23506 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_453
timestamp 0
transform 1 0 23874 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_461
timestamp 0
transform 1 0 24242 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_469
timestamp 0
transform 1 0 24610 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_9_477
timestamp 0
transform 1 0 24978 0 -1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_9_479
timestamp 0
transform 1 0 25070 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_9_481
timestamp 0
transform 1 0 25162 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_489
timestamp 0
transform 1 0 25530 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_497
timestamp 0
transform 1 0 25898 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_9_505
timestamp 0
transform 1 0 26266 0 -1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_9_507
timestamp 0
transform 1 0 26358 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_9_532
timestamp 0
transform 1 0 27508 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_541
timestamp 0
transform 1 0 27922 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_9_573
timestamp 0
transform 1 0 29394 0 -1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_9_581
timestamp 0
transform 1 0 29762 0 -1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_9_585
timestamp 0
transform 1 0 29946 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_10_0
timestamp 0
transform 1 0 3036 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_8
timestamp 0
transform 1 0 3404 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_16
timestamp 0
transform 1 0 3772 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_10_24
timestamp 0
transform 1 0 4140 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_10_28
timestamp 0
transform 1 0 4324 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_10_31
timestamp 0
transform 1 0 4462 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_39
timestamp 0
transform 1 0 4830 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_10_47
timestamp 0
transform 1 0 5198 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_10_51
timestamp 0
transform 1 0 5382 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_10_76
timestamp 0
transform 1 0 6532 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_10_80
timestamp 0
transform 1 0 6716 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_10_86
timestamp 0
transform 1 0 6992 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_10_91
timestamp 0
transform 1 0 7222 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_10_104
timestamp 0
transform 1 0 7820 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_112
timestamp 0
transform 1 0 8188 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_120
timestamp 0
transform 1 0 8556 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_128
timestamp 0
transform 1 0 8924 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_136
timestamp 0
transform 1 0 9292 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_10_144
timestamp 0
transform 1 0 9660 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_10_148
timestamp 0
transform 1 0 9844 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_10_151
timestamp 0
transform 1 0 9982 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_159
timestamp 0
transform 1 0 10350 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_167
timestamp 0
transform 1 0 10718 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_10_175
timestamp 0
transform 1 0 11086 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_10_180
timestamp 0
transform 1 0 11316 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_188
timestamp 0
transform 1 0 11684 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_196
timestamp 0
transform 1 0 12052 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_10_204
timestamp 0
transform 1 0 12420 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_10_208
timestamp 0
transform 1 0 12604 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_10_211
timestamp 0
transform 1 0 12742 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_219
timestamp 0
transform 1 0 13110 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_227
timestamp 0
transform 1 0 13478 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_235
timestamp 0
transform 1 0 13846 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_243
timestamp 0
transform 1 0 14214 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_251
timestamp 0
transform 1 0 14582 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_259
timestamp 0
transform 1 0 14950 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_10_267
timestamp 0
transform 1 0 15318 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_10_269
timestamp 0
transform 1 0 15410 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_10_271
timestamp 0
transform 1 0 15502 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_279
timestamp 0
transform 1 0 15870 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_287
timestamp 0
transform 1 0 16238 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_295
timestamp 0
transform 1 0 16606 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_303
timestamp 0
transform 1 0 16974 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_311
timestamp 0
transform 1 0 17342 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_319
timestamp 0
transform 1 0 17710 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_10_327
timestamp 0
transform 1 0 18078 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_10_329
timestamp 0
transform 1 0 18170 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_10_331
timestamp 0
transform 1 0 18262 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_339
timestamp 0
transform 1 0 18630 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_347
timestamp 0
transform 1 0 18998 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_355
timestamp 0
transform 1 0 19366 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_10_363
timestamp 0
transform 1 0 19734 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_10_365
timestamp 0
transform 1 0 19826 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_10_374
timestamp 0
transform 1 0 20240 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_382
timestamp 0
transform 1 0 20608 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_391
timestamp 0
transform 1 0 21022 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_399
timestamp 0
transform 1 0 21390 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_407
timestamp 0
transform 1 0 21758 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_415
timestamp 0
transform 1 0 22126 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_423
timestamp 0
transform 1 0 22494 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_431
timestamp 0
transform 1 0 22862 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_439
timestamp 0
transform 1 0 23230 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_10_447
timestamp 0
transform 1 0 23598 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_10_449
timestamp 0
transform 1 0 23690 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_10_451
timestamp 0
transform 1 0 23782 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_459
timestamp 0
transform 1 0 24150 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_467
timestamp 0
transform 1 0 24518 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_475
timestamp 0
transform 1 0 24886 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_483
timestamp 0
transform 1 0 25254 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_491
timestamp 0
transform 1 0 25622 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_499
timestamp 0
transform 1 0 25990 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_10_507
timestamp 0
transform 1 0 26358 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_10_509
timestamp 0
transform 1 0 26450 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_10_511
timestamp 0
transform 1 0 26542 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_519
timestamp 0
transform 1 0 26910 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_527
timestamp 0
transform 1 0 27278 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_535
timestamp 0
transform 1 0 27646 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_543
timestamp 0
transform 1 0 28014 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_551
timestamp 0
transform 1 0 28382 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_10_559
timestamp 0
transform 1 0 28750 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_10_567
timestamp 0
transform 1 0 29118 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_10_569
timestamp 0
transform 1 0 29210 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_10_571
timestamp 0
transform 1 0 29302 0 1 5984
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_10_579
timestamp 0
transform 1 0 29670 0 1 5984
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_10_583
timestamp 0
transform 1 0 29854 0 1 5984
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_10_585
timestamp 0
transform 1 0 29946 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_11_0
timestamp 0
transform 1 0 3036 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_8
timestamp 0
transform 1 0 3404 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_16
timestamp 0
transform 1 0 3772 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_24
timestamp 0
transform 1 0 4140 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_32
timestamp 0
transform 1 0 4508 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_40
timestamp 0
transform 1 0 4876 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_48
timestamp 0
transform 1 0 5244 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_11_56
timestamp 0
transform 1 0 5612 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_11_61
timestamp 0
transform 1 0 5842 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_11_72
timestamp 0
transform 1 0 6348 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_11_76
timestamp 0
transform 1 0 6532 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_11_100
timestamp 0
transform 1 0 7636 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_108
timestamp 0
transform 1 0 8004 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_11_116
timestamp 0
transform 1 0 8372 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_11_121
timestamp 0
transform 1 0 8602 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_129
timestamp 0
transform 1 0 8970 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_137
timestamp 0
transform 1 0 9338 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_145
timestamp 0
transform 1 0 9706 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_153
timestamp 0
transform 1 0 10074 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_161
timestamp 0
transform 1 0 10442 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_169
timestamp 0
transform 1 0 10810 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 0
transform 1 0 11178 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_11_179
timestamp 0
transform 1 0 11270 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_11_181
timestamp 0
transform 1 0 11362 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_189
timestamp 0
transform 1 0 11730 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_197
timestamp 0
transform 1 0 12098 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_205
timestamp 0
transform 1 0 12466 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_213
timestamp 0
transform 1 0 12834 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_221
timestamp 0
transform 1 0 13202 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_229
timestamp 0
transform 1 0 13570 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_11_237
timestamp 0
transform 1 0 13938 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_11_239
timestamp 0
transform 1 0 14030 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_11_241
timestamp 0
transform 1 0 14122 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_249
timestamp 0
transform 1 0 14490 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_257
timestamp 0
transform 1 0 14858 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_265
timestamp 0
transform 1 0 15226 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_273
timestamp 0
transform 1 0 15594 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_285
timestamp 0
transform 1 0 16146 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_11_296
timestamp 0
transform 1 0 16652 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_11_301
timestamp 0
transform 1 0 16882 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_11_310
timestamp 0
transform 1 0 17296 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_318
timestamp 0
transform 1 0 17664 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_11_326
timestamp 0
transform 1 0 18032 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_11_337
timestamp 0
transform 1 0 18538 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_11_345
timestamp 0
transform 1 0 18906 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_11_356
timestamp 0
transform 1 0 19412 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_11_361
timestamp 0
transform 1 0 19642 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_11_369
timestamp 0
transform 1 0 20010 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_11_382
timestamp 0
transform 1 0 20608 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 0
transform 1 0 20976 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_11_416
timestamp 0
transform 1 0 22172 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_11_421
timestamp 0
transform 1 0 22402 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_429
timestamp 0
transform 1 0 22770 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_11_461
timestamp 0
transform 1 0 24242 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_11_472
timestamp 0
transform 1 0 24748 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_481
timestamp 0
transform 1 0 25162 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_489
timestamp 0
transform 1 0 25530 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_497
timestamp 0
transform 1 0 25898 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_505
timestamp 0
transform 1 0 26266 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_513
timestamp 0
transform 1 0 26634 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_521
timestamp 0
transform 1 0 27002 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_11_529
timestamp 0
transform 1 0 27370 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_11_537
timestamp 0
transform 1 0 27738 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_11_539
timestamp 0
transform 1 0 27830 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_11_541
timestamp 0
transform 1 0 27922 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_11_545
timestamp 0
transform 1 0 28106 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_11_571
timestamp 0
transform 1 0 29302 0 -1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_11_579
timestamp 0
transform 1 0 29670 0 -1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_11_583
timestamp 0
transform 1 0 29854 0 -1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_11_585
timestamp 0
transform 1 0 29946 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_12_0
timestamp 0
transform 1 0 3036 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_8
timestamp 0
transform 1 0 3404 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_16
timestamp 0
transform 1 0 3772 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_24
timestamp 0
transform 1 0 4140 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_28
timestamp 0
transform 1 0 4324 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_12_31
timestamp 0
transform 1 0 4462 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_39
timestamp 0
transform 1 0 4830 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_47
timestamp 0
transform 1 0 5198 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_55
timestamp 0
transform 1 0 5566 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_67
timestamp 0
transform 1 0 6118 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_75
timestamp 0
transform 1 0 6486 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 0
transform 1 0 6670 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_12_81
timestamp 0
transform 1 0 6762 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_12_86
timestamp 0
transform 1 0 6992 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_12_91
timestamp 0
transform 1 0 7222 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_99
timestamp 0
transform 1 0 7590 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_107
timestamp 0
transform 1 0 7958 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_115
timestamp 0
transform 1 0 8326 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_123
timestamp 0
transform 1 0 8694 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_131
timestamp 0
transform 1 0 9062 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_139
timestamp 0
transform 1 0 9430 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_12_147
timestamp 0
transform 1 0 9798 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_12_149
timestamp 0
transform 1 0 9890 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_12_151
timestamp 0
transform 1 0 9982 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_159
timestamp 0
transform 1 0 10350 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 0
transform 1 0 10718 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_12_192
timestamp 0
transform 1 0 11868 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_200
timestamp 0
transform 1 0 12236 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_12_208
timestamp 0
transform 1 0 12604 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_12_211
timestamp 0
transform 1 0 12742 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_219
timestamp 0
transform 1 0 13110 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_227
timestamp 0
transform 1 0 13478 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_12_231
timestamp 0
transform 1 0 13662 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_12_248
timestamp 0
transform 1 0 14444 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_256
timestamp 0
transform 1 0 14812 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_264
timestamp 0
transform 1 0 15180 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_268
timestamp 0
transform 1 0 15364 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_12_271
timestamp 0
transform 1 0 15502 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_279
timestamp 0
transform 1 0 15870 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_287
timestamp 0
transform 1 0 16238 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_295
timestamp 0
transform 1 0 16606 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_303
timestamp 0
transform 1 0 16974 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_311
timestamp 0
transform 1 0 17342 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_12_319
timestamp 0
transform 1 0 17710 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_12_321
timestamp 0
transform 1 0 17802 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_12_325
timestamp 0
transform 1 0 17986 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_12_329
timestamp 0
transform 1 0 18170 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_12_331
timestamp 0
transform 1 0 18262 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_339
timestamp 0
transform 1 0 18630 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_343
timestamp 0
transform 1 0 18814 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_12_354
timestamp 0
transform 1 0 19320 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_12_358
timestamp 0
transform 1 0 19504 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_12_368
timestamp 0
transform 1 0 19964 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_376
timestamp 0
transform 1 0 20332 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_384
timestamp 0
transform 1 0 20700 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_388
timestamp 0
transform 1 0 20884 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_12_391
timestamp 0
transform 1 0 21022 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_12_419
timestamp 0
transform 1 0 22310 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_427
timestamp 0
transform 1 0 22678 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_435
timestamp 0
transform 1 0 23046 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_443
timestamp 0
transform 1 0 23414 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_447
timestamp 0
transform 1 0 23598 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_12_449
timestamp 0
transform 1 0 23690 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_12_451
timestamp 0
transform 1 0 23782 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_12_479
timestamp 0
transform 1 0 25070 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_487
timestamp 0
transform 1 0 25438 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_495
timestamp 0
transform 1 0 25806 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_503
timestamp 0
transform 1 0 26174 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_507
timestamp 0
transform 1 0 26358 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_12_509
timestamp 0
transform 1 0 26450 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_12_511
timestamp 0
transform 1 0 26542 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_519
timestamp 0
transform 1 0 26910 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_12_527
timestamp 0
transform 1 0 27278 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_535
timestamp 0
transform 1 0 27646 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_539
timestamp 0
transform 1 0 27830 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_12_541
timestamp 0
transform 1 0 27922 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_12_566
timestamp 0
transform 1 0 29072 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_12_571
timestamp 0
transform 1 0 29302 0 1 6528
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_12_579
timestamp 0
transform 1 0 29670 0 1 6528
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_12_583
timestamp 0
transform 1 0 29854 0 1 6528
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_12_585
timestamp 0
transform 1 0 29946 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_13_0
timestamp 0
transform 1 0 3036 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_8
timestamp 0
transform 1 0 3404 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_16
timestamp 0
transform 1 0 3772 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_24
timestamp 0
transform 1 0 4140 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_32
timestamp 0
transform 1 0 4508 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_40
timestamp 0
transform 1 0 4876 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_48
timestamp 0
transform 1 0 5244 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_13_56
timestamp 0
transform 1 0 5612 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_13_61
timestamp 0
transform 1 0 5842 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_13_71
timestamp 0
transform 1 0 6302 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_79
timestamp 0
transform 1 0 6670 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_87
timestamp 0
transform 1 0 7038 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_95
timestamp 0
transform 1 0 7406 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_103
timestamp 0
transform 1 0 7774 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 0
transform 1 0 8142 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_13_116
timestamp 0
transform 1 0 8372 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_13_121
timestamp 0
transform 1 0 8602 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_129
timestamp 0
transform 1 0 8970 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_137
timestamp 0
transform 1 0 9338 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_145
timestamp 0
transform 1 0 9706 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_153
timestamp 0
transform 1 0 10074 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_161
timestamp 0
transform 1 0 10442 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 0
transform 1 0 10810 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_13_171
timestamp 0
transform 1 0 10902 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_13_176
timestamp 0
transform 1 0 11132 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_13_181
timestamp 0
transform 1 0 11362 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_189
timestamp 0
transform 1 0 11730 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_197
timestamp 0
transform 1 0 12098 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_205
timestamp 0
transform 1 0 12466 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_213
timestamp 0
transform 1 0 12834 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_221
timestamp 0
transform 1 0 13202 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_13_229
timestamp 0
transform 1 0 13570 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_13_231
timestamp 0
transform 1 0 13662 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_13_236
timestamp 0
transform 1 0 13892 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_13_241
timestamp 0
transform 1 0 14122 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_13_249
timestamp 0
transform 1 0 14490 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_257
timestamp 0
transform 1 0 14858 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_265
timestamp 0
transform 1 0 15226 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_13_273
timestamp 0
transform 1 0 15594 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_13_282
timestamp 0
transform 1 0 16008 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_13_293
timestamp 0
transform 1 0 16514 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 0
transform 1 0 16698 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_13_299
timestamp 0
transform 1 0 16790 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_13_301
timestamp 0
transform 1 0 16882 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_309
timestamp 0
transform 1 0 17250 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_13_317
timestamp 0
transform 1 0 17618 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_13_321
timestamp 0
transform 1 0 17802 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_13_323
timestamp 0
transform 1 0 17894 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_13_333
timestamp 0
transform 1 0 18354 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_341
timestamp 0
transform 1 0 18722 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_349
timestamp 0
transform 1 0 19090 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_13_357
timestamp 0
transform 1 0 19458 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_13_359
timestamp 0
transform 1 0 19550 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_13_361
timestamp 0
transform 1 0 19642 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_13_369
timestamp 0
transform 1 0 20010 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_13_379
timestamp 0
transform 1 0 20470 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_13_387
timestamp 0
transform 1 0 20838 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 0
transform 1 0 21022 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_13_416
timestamp 0
transform 1 0 22172 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_13_421
timestamp 0
transform 1 0 22402 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_13_433
timestamp 0
transform 1 0 22954 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_13_437
timestamp 0
transform 1 0 23138 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_13_439
timestamp 0
transform 1 0 23230 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_13_464
timestamp 0
transform 1 0 24380 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_13_476
timestamp 0
transform 1 0 24932 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_13_481
timestamp 0
transform 1 0 25162 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_13_489
timestamp 0
transform 1 0 25530 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_13_491
timestamp 0
transform 1 0 25622 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_13_516
timestamp 0
transform 1 0 26772 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_524
timestamp 0
transform 1 0 27140 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_532
timestamp 0
transform 1 0 27508 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_541
timestamp 0
transform 1 0 27922 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_549
timestamp 0
transform 1 0 28290 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_557
timestamp 0
transform 1 0 28658 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_13_572
timestamp 0
transform 1 0 29348 0 -1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_13_580
timestamp 0
transform 1 0 29716 0 -1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_13_584
timestamp 0
transform 1 0 29900 0 -1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_14_0
timestamp 0
transform 1 0 3036 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_8
timestamp 0
transform 1 0 3404 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_16
timestamp 0
transform 1 0 3772 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_24
timestamp 0
transform 1 0 4140 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_14_28
timestamp 0
transform 1 0 4324 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_14_31
timestamp 0
transform 1 0 4462 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_39
timestamp 0
transform 1 0 4830 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_47
timestamp 0
transform 1 0 5198 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_14_51
timestamp 0
transform 1 0 5382 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_14_53
timestamp 0
transform 1 0 5474 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_14_77
timestamp 0
transform 1 0 6578 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_85
timestamp 0
transform 1 0 6946 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 0
transform 1 0 7130 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_14_91
timestamp 0
transform 1 0 7222 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_122
timestamp 0
transform 1 0 8648 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_14_135
timestamp 0
transform 1 0 9246 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_14_139
timestamp 0
transform 1 0 9430 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 0
transform 1 0 9522 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_14_146
timestamp 0
transform 1 0 9752 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_14_151
timestamp 0
transform 1 0 9982 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_159
timestamp 0
transform 1 0 10350 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 0
transform 1 0 10534 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_14_188
timestamp 0
transform 1 0 11684 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_14_198
timestamp 0
transform 1 0 12144 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_206
timestamp 0
transform 1 0 12512 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_14_211
timestamp 0
transform 1 0 12742 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_219
timestamp 0
transform 1 0 13110 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_227
timestamp 0
transform 1 0 13478 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_235
timestamp 0
transform 1 0 13846 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_14_246
timestamp 0
transform 1 0 14352 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_254
timestamp 0
transform 1 0 14720 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_262
timestamp 0
transform 1 0 15088 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_271
timestamp 0
transform 1 0 15502 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_279
timestamp 0
transform 1 0 15870 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_287
timestamp 0
transform 1 0 16238 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_295
timestamp 0
transform 1 0 16606 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_303
timestamp 0
transform 1 0 16974 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_311
timestamp 0
transform 1 0 17342 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_319
timestamp 0
transform 1 0 17710 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_14_327
timestamp 0
transform 1 0 18078 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_14_329
timestamp 0
transform 1 0 18170 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_14_331
timestamp 0
transform 1 0 18262 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_14_335
timestamp 0
transform 1 0 18446 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_14_346
timestamp 0
transform 1 0 18952 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_354
timestamp 0
transform 1 0 19320 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_14_366
timestamp 0
transform 1 0 19872 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_374
timestamp 0
transform 1 0 20240 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_382
timestamp 0
transform 1 0 20608 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_391
timestamp 0
transform 1 0 21022 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_399
timestamp 0
transform 1 0 21390 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_407
timestamp 0
transform 1 0 21758 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_14_415
timestamp 0
transform 1 0 22126 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_14_434
timestamp 0
transform 1 0 23000 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_442
timestamp 0
transform 1 0 23368 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_451
timestamp 0
transform 1 0 23782 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_459
timestamp 0
transform 1 0 24150 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_467
timestamp 0
transform 1 0 24518 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_475
timestamp 0
transform 1 0 24886 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_483
timestamp 0
transform 1 0 25254 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_491
timestamp 0
transform 1 0 25622 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_499
timestamp 0
transform 1 0 25990 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_14_507
timestamp 0
transform 1 0 26358 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_14_509
timestamp 0
transform 1 0 26450 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_14_511
timestamp 0
transform 1 0 26542 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_14_539
timestamp 0
transform 1 0 27830 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_547
timestamp 0
transform 1 0 28198 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_14_555
timestamp 0
transform 1 0 28566 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_563
timestamp 0
transform 1 0 28934 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_14_567
timestamp 0
transform 1 0 29118 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_14_569
timestamp 0
transform 1 0 29210 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_14_571
timestamp 0
transform 1 0 29302 0 1 7072
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_14_579
timestamp 0
transform 1 0 29670 0 1 7072
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_14_583
timestamp 0
transform 1 0 29854 0 1 7072
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_14_585
timestamp 0
transform 1 0 29946 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_15_0
timestamp 0
transform 1 0 3036 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_8
timestamp 0
transform 1 0 3404 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_16
timestamp 0
transform 1 0 3772 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_24
timestamp 0
transform 1 0 4140 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_32
timestamp 0
transform 1 0 4508 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_40
timestamp 0
transform 1 0 4876 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_48
timestamp 0
transform 1 0 5244 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_56
timestamp 0
transform 1 0 5612 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_15_61
timestamp 0
transform 1 0 5842 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_15_69
timestamp 0
transform 1 0 6210 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_77
timestamp 0
transform 1 0 6578 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 0
transform 1 0 6946 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_15_87
timestamp 0
transform 1 0 7038 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_15_94
timestamp 0
transform 1 0 7360 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_102
timestamp 0
transform 1 0 7728 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_15_110
timestamp 0
transform 1 0 8096 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 0
transform 1 0 8464 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_15_121
timestamp 0
transform 1 0 8602 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_129
timestamp 0
transform 1 0 8970 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_15_133
timestamp 0
transform 1 0 9154 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_15_139
timestamp 0
transform 1 0 9430 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_15_146
timestamp 0
transform 1 0 9752 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_154
timestamp 0
transform 1 0 10120 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 0
transform 1 0 10304 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_15_163
timestamp 0
transform 1 0 10534 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_15_176
timestamp 0
transform 1 0 11132 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_15_181
timestamp 0
transform 1 0 11362 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_15_189
timestamp 0
transform 1 0 11730 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_197
timestamp 0
transform 1 0 12098 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_205
timestamp 0
transform 1 0 12466 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_213
timestamp 0
transform 1 0 12834 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_221
timestamp 0
transform 1 0 13202 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_229
timestamp 0
transform 1 0 13570 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_15_237
timestamp 0
transform 1 0 13938 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_15_239
timestamp 0
transform 1 0 14030 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_15_241
timestamp 0
transform 1 0 14122 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_249
timestamp 0
transform 1 0 14490 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_257
timestamp 0
transform 1 0 14858 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_272
timestamp 0
transform 1 0 15548 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_280
timestamp 0
transform 1 0 15916 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_288
timestamp 0
transform 1 0 16284 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_296
timestamp 0
transform 1 0 16652 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_15_301
timestamp 0
transform 1 0 16882 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_309
timestamp 0
transform 1 0 17250 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_317
timestamp 0
transform 1 0 17618 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_325
timestamp 0
transform 1 0 17986 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_15_329
timestamp 0
transform 1 0 18170 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_15_333
timestamp 0
transform 1 0 18354 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_15_341
timestamp 0
transform 1 0 18722 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_15_343
timestamp 0
transform 1 0 18814 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_15_353
timestamp 0
transform 1 0 19274 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_15_357
timestamp 0
transform 1 0 19458 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_15_359
timestamp 0
transform 1 0 19550 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_15_361
timestamp 0
transform 1 0 19642 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_15_369
timestamp 0
transform 1 0 20010 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_15_380
timestamp 0
transform 1 0 20516 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_15_395
timestamp 0
transform 1 0 21206 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_403
timestamp 0
transform 1 0 21574 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_411
timestamp 0
transform 1 0 21942 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_15_419
timestamp 0
transform 1 0 22310 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_15_421
timestamp 0
transform 1 0 22402 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_429
timestamp 0
transform 1 0 22770 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_15_437
timestamp 0
transform 1 0 23138 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_15_439
timestamp 0
transform 1 0 23230 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_15_464
timestamp 0
transform 1 0 24380 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_472
timestamp 0
transform 1 0 24748 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_481
timestamp 0
transform 1 0 25162 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_489
timestamp 0
transform 1 0 25530 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_15_493
timestamp 0
transform 1 0 25714 0 -1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_15_519
timestamp 0
transform 1 0 26910 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_527
timestamp 0
transform 1 0 27278 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_15_535
timestamp 0
transform 1 0 27646 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_15_539
timestamp 0
transform 1 0 27830 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_15_541
timestamp 0
transform 1 0 27922 0 -1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_15_569
timestamp 0
transform 1 0 29210 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_15_577
timestamp 0
transform 1 0 29578 0 -1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_15_585
timestamp 0
transform 1 0 29946 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_16_0
timestamp 0
transform 1 0 3036 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_8
timestamp 0
transform 1 0 3404 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_16
timestamp 0
transform 1 0 3772 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_16_24
timestamp 0
transform 1 0 4140 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_16_28
timestamp 0
transform 1 0 4324 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_16_31
timestamp 0
transform 1 0 4462 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_39
timestamp 0
transform 1 0 4830 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_47
timestamp 0
transform 1 0 5198 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_55
timestamp 0
transform 1 0 5566 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_63
timestamp 0
transform 1 0 5934 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_71
timestamp 0
transform 1 0 6302 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 0
transform 1 0 6670 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_16_81
timestamp 0
transform 1 0 6762 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_16_86
timestamp 0
transform 1 0 6992 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_16_91
timestamp 0
transform 1 0 7222 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_16_102
timestamp 0
transform 1 0 7728 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_110
timestamp 0
transform 1 0 8096 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_16_118
timestamp 0
transform 1 0 8464 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 0
transform 1 0 8648 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_16_126
timestamp 0
transform 1 0 8832 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_134
timestamp 0
transform 1 0 9200 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_142
timestamp 0
transform 1 0 9568 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_151
timestamp 0
transform 1 0 9982 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_16_159
timestamp 0
transform 1 0 10350 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_16_186
timestamp 0
transform 1 0 11592 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_194
timestamp 0
transform 1 0 11960 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_202
timestamp 0
transform 1 0 12328 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_211
timestamp 0
transform 1 0 12742 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_219
timestamp 0
transform 1 0 13110 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_16_227
timestamp 0
transform 1 0 13478 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_16_236
timestamp 0
transform 1 0 13892 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_16_248
timestamp 0
transform 1 0 14444 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_256
timestamp 0
transform 1 0 14812 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_16_264
timestamp 0
transform 1 0 15180 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_16_268
timestamp 0
transform 1 0 15364 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_16_271
timestamp 0
transform 1 0 15502 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_16_282
timestamp 0
transform 1 0 16008 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_290
timestamp 0
transform 1 0 16376 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_298
timestamp 0
transform 1 0 16744 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 0
transform 1 0 17112 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_16_308
timestamp 0
transform 1 0 17204 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_16_316
timestamp 0
transform 1 0 17572 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_16_324
timestamp 0
transform 1 0 17940 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_16_328
timestamp 0
transform 1 0 18124 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_16_331
timestamp 0
transform 1 0 18262 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_339
timestamp 0
transform 1 0 18630 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_16_347
timestamp 0
transform 1 0 18998 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_16_357
timestamp 0
transform 1 0 19458 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_16_365
timestamp 0
transform 1 0 19826 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_16_375
timestamp 0
transform 1 0 20286 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_16_383
timestamp 0
transform 1 0 20654 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_16_387
timestamp 0
transform 1 0 20838 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_16_389
timestamp 0
transform 1 0 20930 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_16_391
timestamp 0
transform 1 0 21022 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_16_404
timestamp 0
transform 1 0 21620 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_16_412
timestamp 0
transform 1 0 21988 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_16_434
timestamp 0
transform 1 0 23000 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_442
timestamp 0
transform 1 0 23368 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_451
timestamp 0
transform 1 0 23782 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_459
timestamp 0
transform 1 0 24150 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_467
timestamp 0
transform 1 0 24518 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_475
timestamp 0
transform 1 0 24886 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_483
timestamp 0
transform 1 0 25254 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_491
timestamp 0
transform 1 0 25622 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_499
timestamp 0
transform 1 0 25990 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_16_507
timestamp 0
transform 1 0 26358 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_16_509
timestamp 0
transform 1 0 26450 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_16_511
timestamp 0
transform 1 0 26542 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_16_523
timestamp 0
transform 1 0 27094 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_16_531
timestamp 0
transform 1 0 27462 0 1 7616
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_16_539
timestamp 0
transform 1 0 27830 0 1 7616
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_16_565
timestamp 0
transform 1 0 29026 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_16_569
timestamp 0
transform 1 0 29210 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_16_571
timestamp 0
transform 1 0 29302 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_16_582
timestamp 0
transform 1 0 29808 0 1 7616
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_17_0
timestamp 0
transform 1 0 3036 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_8
timestamp 0
transform 1 0 3404 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_16
timestamp 0
transform 1 0 3772 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_24
timestamp 0
transform 1 0 4140 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_32
timestamp 0
transform 1 0 4508 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_40
timestamp 0
transform 1 0 4876 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_48
timestamp 0
transform 1 0 5244 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_17_56
timestamp 0
transform 1 0 5612 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_17_61
timestamp 0
transform 1 0 5842 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_17_69
timestamp 0
transform 1 0 6210 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_17_79
timestamp 0
transform 1 0 6670 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_17_106
timestamp 0
transform 1 0 7912 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_17_114
timestamp 0
transform 1 0 8280 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 0
transform 1 0 8464 0 -1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_17_121
timestamp 0
transform 1 0 8602 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_129
timestamp 0
transform 1 0 8970 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_137
timestamp 0
transform 1 0 9338 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_145
timestamp 0
transform 1 0 9706 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_153
timestamp 0
transform 1 0 10074 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_17_161
timestamp 0
transform 1 0 10442 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_17_165
timestamp 0
transform 1 0 10626 0 -1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_17_171
timestamp 0
transform 1 0 10902 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_17_179
timestamp 0
transform 1 0 11270 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_17_181
timestamp 0
transform 1 0 11362 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_189
timestamp 0
transform 1 0 11730 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_197
timestamp 0
transform 1 0 12098 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_205
timestamp 0
transform 1 0 12466 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_213
timestamp 0
transform 1 0 12834 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_221
timestamp 0
transform 1 0 13202 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_229
timestamp 0
transform 1 0 13570 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_17_237
timestamp 0
transform 1 0 13938 0 -1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_17_239
timestamp 0
transform 1 0 14030 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_17_241
timestamp 0
transform 1 0 14122 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_17_251
timestamp 0
transform 1 0 14582 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_17_259
timestamp 0
transform 1 0 14950 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_17_263
timestamp 0
transform 1 0 15134 0 -1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_17_272
timestamp 0
transform 1 0 15548 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_280
timestamp 0
transform 1 0 15916 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_288
timestamp 0
transform 1 0 16284 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_17_296
timestamp 0
transform 1 0 16652 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_17_301
timestamp 0
transform 1 0 16882 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_17_313
timestamp 0
transform 1 0 17434 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_321
timestamp 0
transform 1 0 17802 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_17_329
timestamp 0
transform 1 0 18170 0 -1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_17_331
timestamp 0
transform 1 0 18262 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_17_339
timestamp 0
transform 1 0 18630 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_347
timestamp 0
transform 1 0 18998 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_17_355
timestamp 0
transform 1 0 19366 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_17_359
timestamp 0
transform 1 0 19550 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_17_361
timestamp 0
transform 1 0 19642 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_17_369
timestamp 0
transform 1 0 20010 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_17_381
timestamp 0
transform 1 0 20562 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_17_404
timestamp 0
transform 1 0 21620 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_412
timestamp 0
transform 1 0 21988 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_421
timestamp 0
transform 1 0 22402 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_429
timestamp 0
transform 1 0 22770 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_17_437
timestamp 0
transform 1 0 23138 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_17_462
timestamp 0
transform 1 0 24288 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_17_470
timestamp 0
transform 1 0 24656 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_17_476
timestamp 0
transform 1 0 24932 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_17_481
timestamp 0
transform 1 0 25162 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_489
timestamp 0
transform 1 0 25530 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_497
timestamp 0
transform 1 0 25898 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_505
timestamp 0
transform 1 0 26266 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_513
timestamp 0
transform 1 0 26634 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_521
timestamp 0
transform 1 0 27002 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_529
timestamp 0
transform 1 0 27370 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_17_537
timestamp 0
transform 1 0 27738 0 -1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_17_539
timestamp 0
transform 1 0 27830 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_17_541
timestamp 0
transform 1 0 27922 0 -1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_17_569
timestamp 0
transform 1 0 29210 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_17_577
timestamp 0
transform 1 0 29578 0 -1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_17_585
timestamp 0
transform 1 0 29946 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_0
timestamp 0
transform 1 0 3036 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_8
timestamp 0
transform 1 0 3404 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_16
timestamp 0
transform 1 0 3772 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_18_24
timestamp 0
transform 1 0 4140 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_18_28
timestamp 0
transform 1 0 4324 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_18_31
timestamp 0
transform 1 0 4462 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_39
timestamp 0
transform 1 0 4830 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_47
timestamp 0
transform 1 0 5198 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_18_55
timestamp 0
transform 1 0 5566 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 0
transform 1 0 5658 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_81
timestamp 0
transform 1 0 6762 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 0
transform 1 0 7130 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_91
timestamp 0
transform 1 0 7222 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 0
transform 1 0 7590 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_18_120
timestamp 0
transform 1 0 8556 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_18_130
timestamp 0
transform 1 0 9016 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 0
transform 1 0 9200 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_18_140
timestamp 0
transform 1 0 9476 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_18_148
timestamp 0
transform 1 0 9844 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_18_151
timestamp 0
transform 1 0 9982 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_159
timestamp 0
transform 1 0 10350 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_167
timestamp 0
transform 1 0 10718 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_175
timestamp 0
transform 1 0 11086 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_183
timestamp 0
transform 1 0 11454 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_191
timestamp 0
transform 1 0 11822 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_199
timestamp 0
transform 1 0 12190 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_18_207
timestamp 0
transform 1 0 12558 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_18_209
timestamp 0
transform 1 0 12650 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_211
timestamp 0
transform 1 0 12742 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_219
timestamp 0
transform 1 0 13110 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_227
timestamp 0
transform 1 0 13478 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_235
timestamp 0
transform 1 0 13846 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_243
timestamp 0
transform 1 0 14214 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_251
timestamp 0
transform 1 0 14582 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_259
timestamp 0
transform 1 0 14950 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_18_267
timestamp 0
transform 1 0 15318 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_18_269
timestamp 0
transform 1 0 15410 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_271
timestamp 0
transform 1 0 15502 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_279
timestamp 0
transform 1 0 15870 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_287
timestamp 0
transform 1 0 16238 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_295
timestamp 0
transform 1 0 16606 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_303
timestamp 0
transform 1 0 16974 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_311
timestamp 0
transform 1 0 17342 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_319
timestamp 0
transform 1 0 17710 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_18_327
timestamp 0
transform 1 0 18078 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_18_329
timestamp 0
transform 1 0 18170 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_331
timestamp 0
transform 1 0 18262 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_339
timestamp 0
transform 1 0 18630 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_347
timestamp 0
transform 1 0 18998 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_18_355
timestamp 0
transform 1 0 19366 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_18_359
timestamp 0
transform 1 0 19550 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_368
timestamp 0
transform 1 0 19964 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_376
timestamp 0
transform 1 0 20332 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_18_384
timestamp 0
transform 1 0 20700 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_18_388
timestamp 0
transform 1 0 20884 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_18_391
timestamp 0
transform 1 0 21022 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_399
timestamp 0
transform 1 0 21390 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_407
timestamp 0
transform 1 0 21758 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_435
timestamp 0
transform 1 0 23046 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_18_443
timestamp 0
transform 1 0 23414 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_18_447
timestamp 0
transform 1 0 23598 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_18_449
timestamp 0
transform 1 0 23690 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_451
timestamp 0
transform 1 0 23782 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_18_459
timestamp 0
transform 1 0 24150 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_18_469
timestamp 0
transform 1 0 24610 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_477
timestamp 0
transform 1 0 24978 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_485
timestamp 0
transform 1 0 25346 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_493
timestamp 0
transform 1 0 25714 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_501
timestamp 0
transform 1 0 26082 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_18_509
timestamp 0
transform 1 0 26450 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_511
timestamp 0
transform 1 0 26542 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_519
timestamp 0
transform 1 0 26910 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_527
timestamp 0
transform 1 0 27278 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_535
timestamp 0
transform 1 0 27646 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_543
timestamp 0
transform 1 0 28014 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_551
timestamp 0
transform 1 0 28382 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_18_559
timestamp 0
transform 1 0 28750 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_18_567
timestamp 0
transform 1 0 29118 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_18_569
timestamp 0
transform 1 0 29210 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_18_571
timestamp 0
transform 1 0 29302 0 1 8160
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_18_579
timestamp 0
transform 1 0 29670 0 1 8160
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_18_583
timestamp 0
transform 1 0 29854 0 1 8160
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_18_585
timestamp 0
transform 1 0 29946 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_19_0
timestamp 0
transform 1 0 3036 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_8
timestamp 0
transform 1 0 3404 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_16
timestamp 0
transform 1 0 3772 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_24
timestamp 0
transform 1 0 4140 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_32
timestamp 0
transform 1 0 4508 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_40
timestamp 0
transform 1 0 4876 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_48
timestamp 0
transform 1 0 5244 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_19_56
timestamp 0
transform 1 0 5612 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_19_61
timestamp 0
transform 1 0 5842 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_19_69
timestamp 0
transform 1 0 6210 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_19_96
timestamp 0
transform 1 0 7452 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_19_109
timestamp 0
transform 1 0 8050 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 0
transform 1 0 8418 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 0
transform 1 0 8510 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_19_121
timestamp 0
transform 1 0 8602 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_19_125
timestamp 0
transform 1 0 8786 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_19_127
timestamp 0
transform 1 0 8878 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_19_135
timestamp 0
transform 1 0 9246 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_19_145
timestamp 0
transform 1 0 9706 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_153
timestamp 0
transform 1 0 10074 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_19_167
timestamp 0
transform 1 0 10718 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_19_174
timestamp 0
transform 1 0 11040 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_19_178
timestamp 0
transform 1 0 11224 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_19_181
timestamp 0
transform 1 0 11362 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_189
timestamp 0
transform 1 0 11730 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_197
timestamp 0
transform 1 0 12098 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_205
timestamp 0
transform 1 0 12466 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_213
timestamp 0
transform 1 0 12834 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_221
timestamp 0
transform 1 0 13202 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_229
timestamp 0
transform 1 0 13570 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_19_237
timestamp 0
transform 1 0 13938 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_19_239
timestamp 0
transform 1 0 14030 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_19_241
timestamp 0
transform 1 0 14122 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_249
timestamp 0
transform 1 0 14490 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_257
timestamp 0
transform 1 0 14858 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_265
timestamp 0
transform 1 0 15226 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_273
timestamp 0
transform 1 0 15594 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_281
timestamp 0
transform 1 0 15962 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_289
timestamp 0
transform 1 0 16330 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 0
transform 1 0 16698 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_19_299
timestamp 0
transform 1 0 16790 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_19_301
timestamp 0
transform 1 0 16882 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_19_310
timestamp 0
transform 1 0 17296 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_318
timestamp 0
transform 1 0 17664 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_19_326
timestamp 0
transform 1 0 18032 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_19_335
timestamp 0
transform 1 0 18446 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_343
timestamp 0
transform 1 0 18814 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_351
timestamp 0
transform 1 0 19182 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_19_359
timestamp 0
transform 1 0 19550 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_19_361
timestamp 0
transform 1 0 19642 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_369
timestamp 0
transform 1 0 20010 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_377
timestamp 0
transform 1 0 20378 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_385
timestamp 0
transform 1 0 20746 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 0
transform 1 0 21114 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_19_414
timestamp 0
transform 1 0 22080 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_19_418
timestamp 0
transform 1 0 22264 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_19_421
timestamp 0
transform 1 0 22402 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_19_437
timestamp 0
transform 1 0 23138 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_19_441
timestamp 0
transform 1 0 23322 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_19_466
timestamp 0
transform 1 0 24472 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_19_474
timestamp 0
transform 1 0 24840 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_19_478
timestamp 0
transform 1 0 25024 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_19_481
timestamp 0
transform 1 0 25162 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_19_489
timestamp 0
transform 1 0 25530 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_19_493
timestamp 0
transform 1 0 25714 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_19_519
timestamp 0
transform 1 0 26910 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_527
timestamp 0
transform 1 0 27278 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_19_535
timestamp 0
transform 1 0 27646 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_19_539
timestamp 0
transform 1 0 27830 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_19_541
timestamp 0
transform 1 0 27922 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_549
timestamp 0
transform 1 0 28290 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_19_557
timestamp 0
transform 1 0 28658 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_19_564
timestamp 0
transform 1 0 28980 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_19_572
timestamp 0
transform 1 0 29348 0 -1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_19_580
timestamp 0
transform 1 0 29716 0 -1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_19_584
timestamp 0
transform 1 0 29900 0 -1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_20_0
timestamp 0
transform 1 0 3036 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_8
timestamp 0
transform 1 0 3404 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_16
timestamp 0
transform 1 0 3772 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_24
timestamp 0
transform 1 0 4140 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_20_28
timestamp 0
transform 1 0 4324 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_20_31
timestamp 0
transform 1 0 4462 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_39
timestamp 0
transform 1 0 4830 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_47
timestamp 0
transform 1 0 5198 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_55
timestamp 0
transform 1 0 5566 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_66
timestamp 0
transform 1 0 6072 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_74
timestamp 0
transform 1 0 6440 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_82
timestamp 0
transform 1 0 6808 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_91
timestamp 0
transform 1 0 7222 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_104
timestamp 0
transform 1 0 7820 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_111
timestamp 0
transform 1 0 8142 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_119
timestamp 0
transform 1 0 8510 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_127
timestamp 0
transform 1 0 8878 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_135
timestamp 0
transform 1 0 9246 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_143
timestamp 0
transform 1 0 9614 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 0
transform 1 0 9798 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_20_149
timestamp 0
transform 1 0 9890 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_20_151
timestamp 0
transform 1 0 9982 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_182
timestamp 0
transform 1 0 11408 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_190
timestamp 0
transform 1 0 11776 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_198
timestamp 0
transform 1 0 12144 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_206
timestamp 0
transform 1 0 12512 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_211
timestamp 0
transform 1 0 12742 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_219
timestamp 0
transform 1 0 13110 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_20_223
timestamp 0
transform 1 0 13294 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_20_225
timestamp 0
transform 1 0 13386 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_20_242
timestamp 0
transform 1 0 14168 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_252
timestamp 0
transform 1 0 14628 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_260
timestamp 0
transform 1 0 14996 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_20_268
timestamp 0
transform 1 0 15364 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_20_271
timestamp 0
transform 1 0 15502 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_282
timestamp 0
transform 1 0 16008 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_290
timestamp 0
transform 1 0 16376 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_298
timestamp 0
transform 1 0 16744 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_306
timestamp 0
transform 1 0 17112 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_314
timestamp 0
transform 1 0 17480 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_326
timestamp 0
transform 1 0 18032 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_331
timestamp 0
transform 1 0 18262 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_339
timestamp 0
transform 1 0 18630 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_347
timestamp 0
transform 1 0 18998 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_355
timestamp 0
transform 1 0 19366 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_20_359
timestamp 0
transform 1 0 19550 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_20_361
timestamp 0
transform 1 0 19642 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_20_386
timestamp 0
transform 1 0 20792 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_391
timestamp 0
transform 1 0 21022 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_399
timestamp 0
transform 1 0 21390 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_407
timestamp 0
transform 1 0 21758 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_20_411
timestamp 0
transform 1 0 21942 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_20_432
timestamp 0
transform 1 0 22908 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_440
timestamp 0
transform 1 0 23276 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_20_448
timestamp 0
transform 1 0 23644 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_20_451
timestamp 0
transform 1 0 23782 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_459
timestamp 0
transform 1 0 24150 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_467
timestamp 0
transform 1 0 24518 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_475
timestamp 0
transform 1 0 24886 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_483
timestamp 0
transform 1 0 25254 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_491
timestamp 0
transform 1 0 25622 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_499
timestamp 0
transform 1 0 25990 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_20_507
timestamp 0
transform 1 0 26358 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_20_509
timestamp 0
transform 1 0 26450 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_20_511
timestamp 0
transform 1 0 26542 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_20_539
timestamp 0
transform 1 0 27830 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_547
timestamp 0
transform 1 0 28198 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_20_555
timestamp 0
transform 1 0 28566 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_563
timestamp 0
transform 1 0 28934 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_20_567
timestamp 0
transform 1 0 29118 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_20_569
timestamp 0
transform 1 0 29210 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_20_571
timestamp 0
transform 1 0 29302 0 1 8704
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_20_579
timestamp 0
transform 1 0 29670 0 1 8704
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_20_583
timestamp 0
transform 1 0 29854 0 1 8704
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_20_585
timestamp 0
transform 1 0 29946 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_21_0
timestamp 0
transform 1 0 3036 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_8
timestamp 0
transform 1 0 3404 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_16
timestamp 0
transform 1 0 3772 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_24
timestamp 0
transform 1 0 4140 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_32
timestamp 0
transform 1 0 4508 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_40
timestamp 0
transform 1 0 4876 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_48
timestamp 0
transform 1 0 5244 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_21_56
timestamp 0
transform 1 0 5612 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_21_61
timestamp 0
transform 1 0 5842 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_69
timestamp 0
transform 1 0 6210 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_77
timestamp 0
transform 1 0 6578 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_85
timestamp 0
transform 1 0 6946 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_93
timestamp 0
transform 1 0 7314 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_101
timestamp 0
transform 1 0 7682 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_109
timestamp 0
transform 1 0 8050 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_21_117
timestamp 0
transform 1 0 8418 0 -1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 0
transform 1 0 8510 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_21_121
timestamp 0
transform 1 0 8602 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_129
timestamp 0
transform 1 0 8970 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_137
timestamp 0
transform 1 0 9338 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_145
timestamp 0
transform 1 0 9706 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_153
timestamp 0
transform 1 0 10074 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_161
timestamp 0
transform 1 0 10442 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_169
timestamp 0
transform 1 0 10810 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 0
transform 1 0 11178 0 -1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_21_179
timestamp 0
transform 1 0 11270 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_21_181
timestamp 0
transform 1 0 11362 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_189
timestamp 0
transform 1 0 11730 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_197
timestamp 0
transform 1 0 12098 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_205
timestamp 0
transform 1 0 12466 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_213
timestamp 0
transform 1 0 12834 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_221
timestamp 0
transform 1 0 13202 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_21_229
timestamp 0
transform 1 0 13570 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_21_236
timestamp 0
transform 1 0 13892 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_21_241
timestamp 0
transform 1 0 14122 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 0
transform 1 0 14306 0 -1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_21_247
timestamp 0
transform 1 0 14398 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_21_255
timestamp 0
transform 1 0 14766 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_21_263
timestamp 0
transform 1 0 15134 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_21_271
timestamp 0
transform 1 0 15502 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 0
transform 1 0 15870 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_21_296
timestamp 0
transform 1 0 16652 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_21_301
timestamp 0
transform 1 0 16882 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_21_309
timestamp 0
transform 1 0 17250 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_317
timestamp 0
transform 1 0 17618 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_325
timestamp 0
transform 1 0 17986 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_333
timestamp 0
transform 1 0 18354 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_21_341
timestamp 0
transform 1 0 18722 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_21_356
timestamp 0
transform 1 0 19412 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_21_361
timestamp 0
transform 1 0 19642 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_21_389
timestamp 0
transform 1 0 20930 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_397
timestamp 0
transform 1 0 21298 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_405
timestamp 0
transform 1 0 21666 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_21_413
timestamp 0
transform 1 0 22034 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_21_417
timestamp 0
transform 1 0 22218 0 -1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_21_419
timestamp 0
transform 1 0 22310 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_21_421
timestamp 0
transform 1 0 22402 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_21_445
timestamp 0
transform 1 0 23506 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 0
transform 1 0 23690 0 -1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_21_451
timestamp 0
transform 1 0 23782 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_21_476
timestamp 0
transform 1 0 24932 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_21_481
timestamp 0
transform 1 0 25162 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_21_489
timestamp 0
transform 1 0 25530 0 -1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_21_515
timestamp 0
transform 1 0 26726 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_21_527
timestamp 0
transform 1 0 27278 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_21_535
timestamp 0
transform 1 0 27646 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_21_539
timestamp 0
transform 1 0 27830 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_21_541
timestamp 0
transform 1 0 27922 0 -1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_21_569
timestamp 0
transform 1 0 29210 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_21_577
timestamp 0
transform 1 0 29578 0 -1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_21_585
timestamp 0
transform 1 0 29946 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_0
timestamp 0
transform 1 0 3036 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_8
timestamp 0
transform 1 0 3404 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_16
timestamp 0
transform 1 0 3772 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_22_24
timestamp 0
transform 1 0 4140 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_22_28
timestamp 0
transform 1 0 4324 0 1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_22_31
timestamp 0
transform 1 0 4462 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_39
timestamp 0
transform 1 0 4830 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_47
timestamp 0
transform 1 0 5198 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_55
timestamp 0
transform 1 0 5566 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_63
timestamp 0
transform 1 0 5934 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_71
timestamp 0
transform 1 0 6302 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_79
timestamp 0
transform 1 0 6670 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 0
transform 1 0 7038 0 1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 0
transform 1 0 7130 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_91
timestamp 0
transform 1 0 7222 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_22_99
timestamp 0
transform 1 0 7590 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_123
timestamp 0
transform 1 0 8694 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_131
timestamp 0
transform 1 0 9062 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_139
timestamp 0
transform 1 0 9430 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 0
transform 1 0 9798 0 1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 0
transform 1 0 9890 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_151
timestamp 0
transform 1 0 9982 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_159
timestamp 0
transform 1 0 10350 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_167
timestamp 0
transform 1 0 10718 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_175
timestamp 0
transform 1 0 11086 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_183
timestamp 0
transform 1 0 11454 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_191
timestamp 0
transform 1 0 11822 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_199
timestamp 0
transform 1 0 12190 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_22_207
timestamp 0
transform 1 0 12558 0 1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_22_209
timestamp 0
transform 1 0 12650 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_211
timestamp 0
transform 1 0 12742 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_219
timestamp 0
transform 1 0 13110 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_227
timestamp 0
transform 1 0 13478 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_22_235
timestamp 0
transform 1 0 13846 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_22_255
timestamp 0
transform 1 0 14766 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_22_263
timestamp 0
transform 1 0 15134 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_22_267
timestamp 0
transform 1 0 15318 0 1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_22_269
timestamp 0
transform 1 0 15410 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_22_271
timestamp 0
transform 1 0 15502 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_22_275
timestamp 0
transform 1 0 15686 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_280
timestamp 0
transform 1 0 15916 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_288
timestamp 0
transform 1 0 16284 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_296
timestamp 0
transform 1 0 16652 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_304
timestamp 0
transform 1 0 17020 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_312
timestamp 0
transform 1 0 17388 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_320
timestamp 0
transform 1 0 17756 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_22_328
timestamp 0
transform 1 0 18124 0 1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_22_331
timestamp 0
transform 1 0 18262 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_22_339
timestamp 0
transform 1 0 18630 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_22_343
timestamp 0
transform 1 0 18814 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_364
timestamp 0
transform 1 0 19780 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_372
timestamp 0
transform 1 0 20148 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_22_386
timestamp 0
transform 1 0 20792 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_22_391
timestamp 0
transform 1 0 21022 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_399
timestamp 0
transform 1 0 21390 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_407
timestamp 0
transform 1 0 21758 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_435
timestamp 0
transform 1 0 23046 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_22_443
timestamp 0
transform 1 0 23414 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_22_447
timestamp 0
transform 1 0 23598 0 1 9248
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_22_449
timestamp 0
transform 1 0 23690 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_22_451
timestamp 0
transform 1 0 23782 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_22_479
timestamp 0
transform 1 0 25070 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_22_489
timestamp 0
transform 1 0 25530 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_497
timestamp 0
transform 1 0 25898 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_22_505
timestamp 0
transform 1 0 26266 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_22_509
timestamp 0
transform 1 0 26450 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_511
timestamp 0
transform 1 0 26542 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_22_519
timestamp 0
transform 1 0 26910 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_22_525
timestamp 0
transform 1 0 27186 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_22_533
timestamp 0
transform 1 0 27554 0 1 9248
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_22_541
timestamp 0
transform 1 0 27922 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_22_566
timestamp 0
transform 1 0 29072 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_22_571
timestamp 0
transform 1 0 29302 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_22_581
timestamp 0
transform 1 0 29762 0 1 9248
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_22_585
timestamp 0
transform 1 0 29946 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_23_0
timestamp 0
transform 1 0 3036 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_8
timestamp 0
transform 1 0 3404 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_16
timestamp 0
transform 1 0 3772 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_24
timestamp 0
transform 1 0 4140 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_32
timestamp 0
transform 1 0 4508 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_40
timestamp 0
transform 1 0 4876 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_48
timestamp 0
transform 1 0 5244 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_23_56
timestamp 0
transform 1 0 5612 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_23_61
timestamp 0
transform 1 0 5842 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_69
timestamp 0
transform 1 0 6210 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_77
timestamp 0
transform 1 0 6578 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_85
timestamp 0
transform 1 0 6946 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_93
timestamp 0
transform 1 0 7314 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 0
transform 1 0 7682 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_23_103
timestamp 0
transform 1 0 7774 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_23_111
timestamp 0
transform 1 0 8142 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 0
transform 1 0 8510 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_23_121
timestamp 0
transform 1 0 8602 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_23_130
timestamp 0
transform 1 0 9016 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 0
transform 1 0 9384 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_23_145
timestamp 0
transform 1 0 9706 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_23_156
timestamp 0
transform 1 0 10212 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_164
timestamp 0
transform 1 0 10580 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_172
timestamp 0
transform 1 0 10948 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_181
timestamp 0
transform 1 0 11362 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_189
timestamp 0
transform 1 0 11730 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_197
timestamp 0
transform 1 0 12098 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_205
timestamp 0
transform 1 0 12466 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_213
timestamp 0
transform 1 0 12834 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_221
timestamp 0
transform 1 0 13202 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_229
timestamp 0
transform 1 0 13570 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_237
timestamp 0
transform 1 0 13938 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_23_239
timestamp 0
transform 1 0 14030 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_23_241
timestamp 0
transform 1 0 14122 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_23_245
timestamp 0
transform 1 0 14306 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_23_250
timestamp 0
transform 1 0 14536 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_258
timestamp 0
transform 1 0 14904 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_266
timestamp 0
transform 1 0 15272 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_274
timestamp 0
transform 1 0 15640 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_282
timestamp 0
transform 1 0 16008 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_290
timestamp 0
transform 1 0 16376 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_298
timestamp 0
transform 1 0 16744 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_23_301
timestamp 0
transform 1 0 16882 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_23_310
timestamp 0
transform 1 0 17296 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_318
timestamp 0
transform 1 0 17664 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_326
timestamp 0
transform 1 0 18032 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_334
timestamp 0
transform 1 0 18400 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_23_342
timestamp 0
transform 1 0 18768 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_23_346
timestamp 0
transform 1 0 18952 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_23_356
timestamp 0
transform 1 0 19412 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_23_361
timestamp 0
transform 1 0 19642 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_369
timestamp 0
transform 1 0 20010 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_377
timestamp 0
transform 1 0 20378 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_23_379
timestamp 0
transform 1 0 20470 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_23_385
timestamp 0
transform 1 0 20746 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_393
timestamp 0
transform 1 0 21114 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_401
timestamp 0
transform 1 0 21482 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_409
timestamp 0
transform 1 0 21850 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_417
timestamp 0
transform 1 0 22218 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_23_419
timestamp 0
transform 1 0 22310 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_23_421
timestamp 0
transform 1 0 22402 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_23_445
timestamp 0
transform 1 0 23506 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_453
timestamp 0
transform 1 0 23874 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_461
timestamp 0
transform 1 0 24242 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_469
timestamp 0
transform 1 0 24610 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_477
timestamp 0
transform 1 0 24978 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_23_479
timestamp 0
transform 1 0 25070 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_23_481
timestamp 0
transform 1 0 25162 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_489
timestamp 0
transform 1 0 25530 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_497
timestamp 0
transform 1 0 25898 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_505
timestamp 0
transform 1 0 26266 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_513
timestamp 0
transform 1 0 26634 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_521
timestamp 0
transform 1 0 27002 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_529
timestamp 0
transform 1 0 27370 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_23_537
timestamp 0
transform 1 0 27738 0 -1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_23_539
timestamp 0
transform 1 0 27830 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_23_541
timestamp 0
transform 1 0 27922 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_549
timestamp 0
transform 1 0 28290 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_557
timestamp 0
transform 1 0 28658 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_565
timestamp 0
transform 1 0 29026 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_23_573
timestamp 0
transform 1 0 29394 0 -1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_23_581
timestamp 0
transform 1 0 29762 0 -1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_23_585
timestamp 0
transform 1 0 29946 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_24_0
timestamp 0
transform 1 0 3036 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_8
timestamp 0
transform 1 0 3404 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_16
timestamp 0
transform 1 0 3772 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_24_24
timestamp 0
transform 1 0 4140 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_24_28
timestamp 0
transform 1 0 4324 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_24_31
timestamp 0
transform 1 0 4462 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_39
timestamp 0
transform 1 0 4830 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_47
timestamp 0
transform 1 0 5198 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_55
timestamp 0
transform 1 0 5566 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_63
timestamp 0
transform 1 0 5934 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_71
timestamp 0
transform 1 0 6302 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_79
timestamp 0
transform 1 0 6670 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 0
transform 1 0 7038 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_89
timestamp 0
transform 1 0 7130 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_24_91
timestamp 0
transform 1 0 7222 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_24_95
timestamp 0
transform 1 0 7406 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_24_99
timestamp 0
transform 1 0 7590 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_24_126
timestamp 0
transform 1 0 8832 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_24_135
timestamp 0
transform 1 0 9246 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_24_146
timestamp 0
transform 1 0 9752 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_24_151
timestamp 0
transform 1 0 9982 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_24_175
timestamp 0
transform 1 0 11086 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_183
timestamp 0
transform 1 0 11454 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_191
timestamp 0
transform 1 0 11822 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_199
timestamp 0
transform 1 0 12190 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_24_207
timestamp 0
transform 1 0 12558 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_209
timestamp 0
transform 1 0 12650 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_24_211
timestamp 0
transform 1 0 12742 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_219
timestamp 0
transform 1 0 13110 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_227
timestamp 0
transform 1 0 13478 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_235
timestamp 0
transform 1 0 13846 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_24_243
timestamp 0
transform 1 0 14214 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_245
timestamp 0
transform 1 0 14306 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_24_250
timestamp 0
transform 1 0 14536 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_258
timestamp 0
transform 1 0 14904 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_24_266
timestamp 0
transform 1 0 15272 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_24_271
timestamp 0
transform 1 0 15502 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_279
timestamp 0
transform 1 0 15870 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_287
timestamp 0
transform 1 0 16238 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_295
timestamp 0
transform 1 0 16606 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_24_303
timestamp 0
transform 1 0 16974 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_305
timestamp 0
transform 1 0 17066 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_24_315
timestamp 0
transform 1 0 17526 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_24_319
timestamp 0
transform 1 0 17710 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_321
timestamp 0
transform 1 0 17802 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_24_326
timestamp 0
transform 1 0 18032 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_24_331
timestamp 0
transform 1 0 18262 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_24_351
timestamp 0
transform 1 0 19182 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_359
timestamp 0
transform 1 0 19550 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_367
timestamp 0
transform 1 0 19918 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_375
timestamp 0
transform 1 0 20286 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_24_383
timestamp 0
transform 1 0 20654 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_24_387
timestamp 0
transform 1 0 20838 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_389
timestamp 0
transform 1 0 20930 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_24_391
timestamp 0
transform 1 0 21022 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_399
timestamp 0
transform 1 0 21390 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_407
timestamp 0
transform 1 0 21758 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_24_415
timestamp 0
transform 1 0 22126 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_24_428
timestamp 0
transform 1 0 22724 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_436
timestamp 0
transform 1 0 23092 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_24_444
timestamp 0
transform 1 0 23460 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_24_448
timestamp 0
transform 1 0 23644 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_24_451
timestamp 0
transform 1 0 23782 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_459
timestamp 0
transform 1 0 24150 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_467
timestamp 0
transform 1 0 24518 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_475
timestamp 0
transform 1 0 24886 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_483
timestamp 0
transform 1 0 25254 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_491
timestamp 0
transform 1 0 25622 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_499
timestamp 0
transform 1 0 25990 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_24_507
timestamp 0
transform 1 0 26358 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_509
timestamp 0
transform 1 0 26450 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_24_511
timestamp 0
transform 1 0 26542 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_519
timestamp 0
transform 1 0 26910 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_527
timestamp 0
transform 1 0 27278 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_535
timestamp 0
transform 1 0 27646 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_543
timestamp 0
transform 1 0 28014 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_551
timestamp 0
transform 1 0 28382 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_24_559
timestamp 0
transform 1 0 28750 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_24_567
timestamp 0
transform 1 0 29118 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_569
timestamp 0
transform 1 0 29210 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_24_571
timestamp 0
transform 1 0 29302 0 1 9792
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_24_579
timestamp 0
transform 1 0 29670 0 1 9792
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_24_583
timestamp 0
transform 1 0 29854 0 1 9792
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_24_585
timestamp 0
transform 1 0 29946 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_25_0
timestamp 0
transform 1 0 3036 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_8
timestamp 0
transform 1 0 3404 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_16
timestamp 0
transform 1 0 3772 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_24
timestamp 0
transform 1 0 4140 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_32
timestamp 0
transform 1 0 4508 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_40
timestamp 0
transform 1 0 4876 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_48
timestamp 0
transform 1 0 5244 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_25_56
timestamp 0
transform 1 0 5612 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_25_61
timestamp 0
transform 1 0 5842 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_69
timestamp 0
transform 1 0 6210 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_77
timestamp 0
transform 1 0 6578 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_85
timestamp 0
transform 1 0 6946 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_93
timestamp 0
transform 1 0 7314 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_25_101
timestamp 0
transform 1 0 7682 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 0
transform 1 0 7866 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_25_114
timestamp 0
transform 1 0 8280 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 0
transform 1 0 8464 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_25_121
timestamp 0
transform 1 0 8602 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_25_125
timestamp 0
transform 1 0 8786 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_25_131
timestamp 0
transform 1 0 9062 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 0
transform 1 0 9430 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_25_164
timestamp 0
transform 1 0 10580 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_172
timestamp 0
transform 1 0 10948 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_181
timestamp 0
transform 1 0 11362 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_189
timestamp 0
transform 1 0 11730 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_197
timestamp 0
transform 1 0 12098 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_205
timestamp 0
transform 1 0 12466 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_213
timestamp 0
transform 1 0 12834 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_221
timestamp 0
transform 1 0 13202 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_229
timestamp 0
transform 1 0 13570 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_25_237
timestamp 0
transform 1 0 13938 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_25_239
timestamp 0
transform 1 0 14030 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_25_241
timestamp 0
transform 1 0 14122 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_25_261
timestamp 0
transform 1 0 15042 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_25_269
timestamp 0
transform 1 0 15410 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_25_296
timestamp 0
transform 1 0 16652 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_25_301
timestamp 0
transform 1 0 16882 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_309
timestamp 0
transform 1 0 17250 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_317
timestamp 0
transform 1 0 17618 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_325
timestamp 0
transform 1 0 17986 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_333
timestamp 0
transform 1 0 18354 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_341
timestamp 0
transform 1 0 18722 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_349
timestamp 0
transform 1 0 19090 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_25_357
timestamp 0
transform 1 0 19458 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_25_359
timestamp 0
transform 1 0 19550 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_25_361
timestamp 0
transform 1 0 19642 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_369
timestamp 0
transform 1 0 20010 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_377
timestamp 0
transform 1 0 20378 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_385
timestamp 0
transform 1 0 20746 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_393
timestamp 0
transform 1 0 21114 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_401
timestamp 0
transform 1 0 21482 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_409
timestamp 0
transform 1 0 21850 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_25_417
timestamp 0
transform 1 0 22218 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_25_419
timestamp 0
transform 1 0 22310 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_25_421
timestamp 0
transform 1 0 22402 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_429
timestamp 0
transform 1 0 22770 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_437
timestamp 0
transform 1 0 23138 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_445
timestamp 0
transform 1 0 23506 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_453
timestamp 0
transform 1 0 23874 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_461
timestamp 0
transform 1 0 24242 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_469
timestamp 0
transform 1 0 24610 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_25_477
timestamp 0
transform 1 0 24978 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_25_479
timestamp 0
transform 1 0 25070 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_25_481
timestamp 0
transform 1 0 25162 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_25_509
timestamp 0
transform 1 0 26450 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_517
timestamp 0
transform 1 0 26818 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_525
timestamp 0
transform 1 0 27186 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_25_533
timestamp 0
transform 1 0 27554 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_25_537
timestamp 0
transform 1 0 27738 0 -1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_25_539
timestamp 0
transform 1 0 27830 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_25_541
timestamp 0
transform 1 0 27922 0 -1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_25_569
timestamp 0
transform 1 0 29210 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_25_577
timestamp 0
transform 1 0 29578 0 -1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_25_585
timestamp 0
transform 1 0 29946 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_0
timestamp 0
transform 1 0 3036 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_8
timestamp 0
transform 1 0 3404 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_16
timestamp 0
transform 1 0 3772 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_26_24
timestamp 0
transform 1 0 4140 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_26_28
timestamp 0
transform 1 0 4324 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_26_31
timestamp 0
transform 1 0 4462 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_26_39
timestamp 0
transform 1 0 4830 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_26_41
timestamp 0
transform 1 0 4922 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_65
timestamp 0
transform 1 0 6026 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_73
timestamp 0
transform 1 0 6394 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_81
timestamp 0
transform 1 0 6762 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 0
transform 1 0 7130 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_91
timestamp 0
transform 1 0 7222 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_99
timestamp 0
transform 1 0 7590 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_107
timestamp 0
transform 1 0 7958 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_26_120
timestamp 0
transform 1 0 8556 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_26_144
timestamp 0
transform 1 0 9660 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_26_148
timestamp 0
transform 1 0 9844 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_26_151
timestamp 0
transform 1 0 9982 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_159
timestamp 0
transform 1 0 10350 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_167
timestamp 0
transform 1 0 10718 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_175
timestamp 0
transform 1 0 11086 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_183
timestamp 0
transform 1 0 11454 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_191
timestamp 0
transform 1 0 11822 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_199
timestamp 0
transform 1 0 12190 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_26_207
timestamp 0
transform 1 0 12558 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_26_209
timestamp 0
transform 1 0 12650 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_211
timestamp 0
transform 1 0 12742 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_219
timestamp 0
transform 1 0 13110 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_26_227
timestamp 0
transform 1 0 13478 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_26_251
timestamp 0
transform 1 0 14582 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_26_259
timestamp 0
transform 1 0 14950 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_26_267
timestamp 0
transform 1 0 15318 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_26_269
timestamp 0
transform 1 0 15410 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_271
timestamp 0
transform 1 0 15502 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_26_302
timestamp 0
transform 1 0 16928 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_26_315
timestamp 0
transform 1 0 17526 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_26_323
timestamp 0
transform 1 0 17894 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_26_327
timestamp 0
transform 1 0 18078 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_26_329
timestamp 0
transform 1 0 18170 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_331
timestamp 0
transform 1 0 18262 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_342
timestamp 0
transform 1 0 18768 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_26_350
timestamp 0
transform 1 0 19136 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_26_354
timestamp 0
transform 1 0 19320 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_379
timestamp 0
transform 1 0 20470 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_26_387
timestamp 0
transform 1 0 20838 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_26_389
timestamp 0
transform 1 0 20930 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_391
timestamp 0
transform 1 0 21022 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_399
timestamp 0
transform 1 0 21390 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_407
timestamp 0
transform 1 0 21758 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_415
timestamp 0
transform 1 0 22126 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_423
timestamp 0
transform 1 0 22494 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_26_431
timestamp 0
transform 1 0 22862 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_26_433
timestamp 0
transform 1 0 22954 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_26_437
timestamp 0
transform 1 0 23138 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_26_445
timestamp 0
transform 1 0 23506 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_26_449
timestamp 0
transform 1 0 23690 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_26_451
timestamp 0
transform 1 0 23782 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_26_459
timestamp 0
transform 1 0 24150 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_26_467
timestamp 0
transform 1 0 24518 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_26_493
timestamp 0
transform 1 0 25714 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_26_505
timestamp 0
transform 1 0 26266 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_26_509
timestamp 0
transform 1 0 26450 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_26_511
timestamp 0
transform 1 0 26542 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_26_519
timestamp 0
transform 1 0 26910 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_26_527
timestamp 0
transform 1 0 27278 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 0
transform 1 0 27462 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_26_556
timestamp 0
transform 1 0 28612 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_26_566
timestamp 0
transform 1 0 29072 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_26_571
timestamp 0
transform 1 0 29302 0 1 10336
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_26_579
timestamp 0
transform 1 0 29670 0 1 10336
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_26_583
timestamp 0
transform 1 0 29854 0 1 10336
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_26_585
timestamp 0
transform 1 0 29946 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_27_0
timestamp 0
transform 1 0 3036 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_8
timestamp 0
transform 1 0 3404 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_16
timestamp 0
transform 1 0 3772 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_24
timestamp 0
transform 1 0 4140 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_32
timestamp 0
transform 1 0 4508 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_40
timestamp 0
transform 1 0 4876 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_48
timestamp 0
transform 1 0 5244 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_56
timestamp 0
transform 1 0 5612 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_27_61
timestamp 0
transform 1 0 5842 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_69
timestamp 0
transform 1 0 6210 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_77
timestamp 0
transform 1 0 6578 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_85
timestamp 0
transform 1 0 6946 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_93
timestamp 0
transform 1 0 7314 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_101
timestamp 0
transform 1 0 7682 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_109
timestamp 0
transform 1 0 8050 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_27_117
timestamp 0
transform 1 0 8418 0 -1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 0
transform 1 0 8510 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_27_121
timestamp 0
transform 1 0 8602 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_129
timestamp 0
transform 1 0 8970 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_137
timestamp 0
transform 1 0 9338 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_145
timestamp 0
transform 1 0 9706 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 0
transform 1 0 9890 0 -1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 0
transform 1 0 9982 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_27_176
timestamp 0
transform 1 0 11132 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_27_181
timestamp 0
transform 1 0 11362 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_27_185
timestamp 0
transform 1 0 11546 0 -1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_27_187
timestamp 0
transform 1 0 11638 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_27_199
timestamp 0
transform 1 0 12190 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_27_227
timestamp 0
transform 1 0 13478 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_235
timestamp 0
transform 1 0 13846 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_27_239
timestamp 0
transform 1 0 14030 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_27_241
timestamp 0
transform 1 0 14122 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_27_245
timestamp 0
transform 1 0 14306 0 -1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 0
transform 1 0 14398 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_27_272
timestamp 0
transform 1 0 15548 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_27_287
timestamp 0
transform 1 0 16238 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_295
timestamp 0
transform 1 0 16606 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_27_299
timestamp 0
transform 1 0 16790 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_27_301
timestamp 0
transform 1 0 16882 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_309
timestamp 0
transform 1 0 17250 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_317
timestamp 0
transform 1 0 17618 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_325
timestamp 0
transform 1 0 17986 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_27_336
timestamp 0
transform 1 0 18492 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_27_356
timestamp 0
transform 1 0 19412 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_27_361
timestamp 0
transform 1 0 19642 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_369
timestamp 0
transform 1 0 20010 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_27_377
timestamp 0
transform 1 0 20378 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_385
timestamp 0
transform 1 0 20746 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_27_389
timestamp 0
transform 1 0 20930 0 -1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 0
transform 1 0 21022 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_27_416
timestamp 0
transform 1 0 22172 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_27_421
timestamp 0
transform 1 0 22402 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_27_429
timestamp 0
transform 1 0 22770 0 -1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_27_431
timestamp 0
transform 1 0 22862 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_27_435
timestamp 0
transform 1 0 23046 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_27_455
timestamp 0
transform 1 0 23966 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_27_475
timestamp 0
transform 1 0 24886 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_27_479
timestamp 0
transform 1 0 25070 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_27_481
timestamp 0
transform 1 0 25162 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_27_509
timestamp 0
transform 1 0 26450 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_27_513
timestamp 0
transform 1 0 26634 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_27_518
timestamp 0
transform 1 0 26864 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_526
timestamp 0
transform 1 0 27232 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_27_534
timestamp 0
transform 1 0 27600 0 -1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_27_538
timestamp 0
transform 1 0 27784 0 -1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_27_541
timestamp 0
transform 1 0 27922 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_549
timestamp 0
transform 1 0 28290 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_557
timestamp 0
transform 1 0 28658 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_569
timestamp 0
transform 1 0 29210 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_27_577
timestamp 0
transform 1 0 29578 0 -1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_27_585
timestamp 0
transform 1 0 29946 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_28_0
timestamp 0
transform 1 0 3036 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_8
timestamp 0
transform 1 0 3404 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_16
timestamp 0
transform 1 0 3772 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_28_24
timestamp 0
transform 1 0 4140 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_28_28
timestamp 0
transform 1 0 4324 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_28_31
timestamp 0
transform 1 0 4462 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_28_39
timestamp 0
transform 1 0 4830 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_28_52
timestamp 0
transform 1 0 5428 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_28_80
timestamp 0
transform 1 0 6716 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 0
transform 1 0 7084 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_28_91
timestamp 0
transform 1 0 7222 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_99
timestamp 0
transform 1 0 7590 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_107
timestamp 0
transform 1 0 7958 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_115
timestamp 0
transform 1 0 8326 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_123
timestamp 0
transform 1 0 8694 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_131
timestamp 0
transform 1 0 9062 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_139
timestamp 0
transform 1 0 9430 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 0
transform 1 0 9798 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_28_149
timestamp 0
transform 1 0 9890 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_28_151
timestamp 0
transform 1 0 9982 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_159
timestamp 0
transform 1 0 10350 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_28_167
timestamp 0
transform 1 0 10718 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_28_193
timestamp 0
transform 1 0 11914 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_201
timestamp 0
transform 1 0 12282 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_28_209
timestamp 0
transform 1 0 12650 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_28_211
timestamp 0
transform 1 0 12742 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_219
timestamp 0
transform 1 0 13110 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_28_227
timestamp 0
transform 1 0 13478 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_28_240
timestamp 0
transform 1 0 14076 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_248
timestamp 0
transform 1 0 14444 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_256
timestamp 0
transform 1 0 14812 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_28_264
timestamp 0
transform 1 0 15180 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_28_268
timestamp 0
transform 1 0 15364 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_28_271
timestamp 0
transform 1 0 15502 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_28_279
timestamp 0
transform 1 0 15870 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_28_283
timestamp 0
transform 1 0 16054 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_28_291
timestamp 0
transform 1 0 16422 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_312
timestamp 0
transform 1 0 17388 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_320
timestamp 0
transform 1 0 17756 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_28_328
timestamp 0
transform 1 0 18124 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_28_331
timestamp 0
transform 1 0 18262 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_28_339
timestamp 0
transform 1 0 18630 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_347
timestamp 0
transform 1 0 18998 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_355
timestamp 0
transform 1 0 19366 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_363
timestamp 0
transform 1 0 19734 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_371
timestamp 0
transform 1 0 20102 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_379
timestamp 0
transform 1 0 20470 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_28_387
timestamp 0
transform 1 0 20838 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_28_389
timestamp 0
transform 1 0 20930 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_28_391
timestamp 0
transform 1 0 21022 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_28_419
timestamp 0
transform 1 0 22310 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_28_429
timestamp 0
transform 1 0 22770 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_440
timestamp 0
transform 1 0 23276 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_28_448
timestamp 0
transform 1 0 23644 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_28_451
timestamp 0
transform 1 0 23782 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_28_458
timestamp 0
transform 1 0 24104 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_466
timestamp 0
transform 1 0 24472 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_474
timestamp 0
transform 1 0 24840 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_482
timestamp 0
transform 1 0 25208 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_490
timestamp 0
transform 1 0 25576 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_498
timestamp 0
transform 1 0 25944 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_28_506
timestamp 0
transform 1 0 26312 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_28_511
timestamp 0
transform 1 0 26542 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_519
timestamp 0
transform 1 0 26910 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_527
timestamp 0
transform 1 0 27278 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_535
timestamp 0
transform 1 0 27646 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_543
timestamp 0
transform 1 0 28014 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_551
timestamp 0
transform 1 0 28382 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_28_559
timestamp 0
transform 1 0 28750 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_28_567
timestamp 0
transform 1 0 29118 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_28_569
timestamp 0
transform 1 0 29210 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_28_571
timestamp 0
transform 1 0 29302 0 1 10880
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_28_579
timestamp 0
transform 1 0 29670 0 1 10880
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_28_583
timestamp 0
transform 1 0 29854 0 1 10880
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_28_585
timestamp 0
transform 1 0 29946 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_29_0
timestamp 0
transform 1 0 3036 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_8
timestamp 0
transform 1 0 3404 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_16
timestamp 0
transform 1 0 3772 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_24
timestamp 0
transform 1 0 4140 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_29_56
timestamp 0
transform 1 0 5612 0 -1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_29_61
timestamp 0
transform 1 0 5842 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_69
timestamp 0
transform 1 0 6210 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_101
timestamp 0
transform 1 0 7682 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_109
timestamp 0
transform 1 0 8050 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_117
timestamp 0
transform 1 0 8418 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 0
transform 1 0 8510 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_29_121
timestamp 0
transform 1 0 8602 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_129
timestamp 0
transform 1 0 8970 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_137
timestamp 0
transform 1 0 9338 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_145
timestamp 0
transform 1 0 9706 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_153
timestamp 0
transform 1 0 10074 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_161
timestamp 0
transform 1 0 10442 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_169
timestamp 0
transform 1 0 10810 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_177
timestamp 0
transform 1 0 11178 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_29_179
timestamp 0
transform 1 0 11270 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_29_181
timestamp 0
transform 1 0 11362 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_189
timestamp 0
transform 1 0 11730 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_197
timestamp 0
transform 1 0 12098 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_205
timestamp 0
transform 1 0 12466 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_213
timestamp 0
transform 1 0 12834 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_221
timestamp 0
transform 1 0 13202 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_229
timestamp 0
transform 1 0 13570 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 0
transform 1 0 13938 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_29_239
timestamp 0
transform 1 0 14030 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_29_241
timestamp 0
transform 1 0 14122 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_249
timestamp 0
transform 1 0 14490 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_257
timestamp 0
transform 1 0 14858 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_265
timestamp 0
transform 1 0 15226 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_273
timestamp 0
transform 1 0 15594 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 0
transform 1 0 15962 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_29_289
timestamp 0
transform 1 0 16330 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_297
timestamp 0
transform 1 0 16698 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_29_299
timestamp 0
transform 1 0 16790 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_29_301
timestamp 0
transform 1 0 16882 0 -1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_29_309
timestamp 0
transform 1 0 17250 0 -1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_29_316
timestamp 0
transform 1 0 17572 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_324
timestamp 0
transform 1 0 17940 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_332
timestamp 0
transform 1 0 18308 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_29_334
timestamp 0
transform 1 0 18400 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_29_338
timestamp 0
transform 1 0 18584 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_346
timestamp 0
transform 1 0 18952 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_29_354
timestamp 0
transform 1 0 19320 0 -1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_29_358
timestamp 0
transform 1 0 19504 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_29_361
timestamp 0
transform 1 0 19642 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_369
timestamp 0
transform 1 0 20010 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_377
timestamp 0
transform 1 0 20378 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_29_403
timestamp 0
transform 1 0 21574 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_411
timestamp 0
transform 1 0 21942 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_29_419
timestamp 0
transform 1 0 22310 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_29_421
timestamp 0
transform 1 0 22402 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_429
timestamp 0
transform 1 0 22770 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_437
timestamp 0
transform 1 0 23138 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_445
timestamp 0
transform 1 0 23506 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_453
timestamp 0
transform 1 0 23874 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_461
timestamp 0
transform 1 0 24242 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_29_469
timestamp 0
transform 1 0 24610 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_477
timestamp 0
transform 1 0 24978 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_29_479
timestamp 0
transform 1 0 25070 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_29_481
timestamp 0
transform 1 0 25162 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_489
timestamp 0
transform 1 0 25530 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_497
timestamp 0
transform 1 0 25898 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_505
timestamp 0
transform 1 0 26266 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_513
timestamp 0
transform 1 0 26634 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_521
timestamp 0
transform 1 0 27002 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_29_529
timestamp 0
transform 1 0 27370 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_537
timestamp 0
transform 1 0 27738 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_29_539
timestamp 0
transform 1 0 27830 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_29_541
timestamp 0
transform 1 0 27922 0 -1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_29_569
timestamp 0
transform 1 0 29210 0 -1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_29_576
timestamp 0
transform 1 0 29532 0 -1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_29_584
timestamp 0
transform 1 0 29900 0 -1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_30_0
timestamp 0
transform 1 0 3036 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_8
timestamp 0
transform 1 0 3404 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_16
timestamp 0
transform 1 0 3772 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_24
timestamp 0
transform 1 0 4140 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_30_28
timestamp 0
transform 1 0 4324 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_30_31
timestamp 0
transform 1 0 4462 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_39
timestamp 0
transform 1 0 4830 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_47
timestamp 0
transform 1 0 5198 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_55
timestamp 0
transform 1 0 5566 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 0
transform 1 0 5750 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 0
transform 1 0 5842 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_30_86
timestamp 0
transform 1 0 6992 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_30_91
timestamp 0
transform 1 0 7222 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_30_102
timestamp 0
transform 1 0 7728 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_110
timestamp 0
transform 1 0 8096 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_118
timestamp 0
transform 1 0 8464 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_30_146
timestamp 0
transform 1 0 9752 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_30_151
timestamp 0
transform 1 0 9982 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_30_159
timestamp 0
transform 1 0 10350 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_167
timestamp 0
transform 1 0 10718 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 0
transform 1 0 10902 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_30_196
timestamp 0
transform 1 0 12052 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_204
timestamp 0
transform 1 0 12420 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_30_208
timestamp 0
transform 1 0 12604 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_30_211
timestamp 0
transform 1 0 12742 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_30_239
timestamp 0
transform 1 0 14030 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_247
timestamp 0
transform 1 0 14398 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_255
timestamp 0
transform 1 0 14766 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_263
timestamp 0
transform 1 0 15134 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_30_267
timestamp 0
transform 1 0 15318 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_30_269
timestamp 0
transform 1 0 15410 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_30_271
timestamp 0
transform 1 0 15502 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_279
timestamp 0
transform 1 0 15870 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_30_287
timestamp 0
transform 1 0 16238 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_30_293
timestamp 0
transform 1 0 16514 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_301
timestamp 0
transform 1 0 16882 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_309
timestamp 0
transform 1 0 17250 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_317
timestamp 0
transform 1 0 17618 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_325
timestamp 0
transform 1 0 17986 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_30_329
timestamp 0
transform 1 0 18170 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_30_331
timestamp 0
transform 1 0 18262 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_342
timestamp 0
transform 1 0 18768 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_350
timestamp 0
transform 1 0 19136 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_30_354
timestamp 0
transform 1 0 19320 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_30_361
timestamp 0
transform 1 0 19642 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_369
timestamp 0
transform 1 0 20010 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_377
timestamp 0
transform 1 0 20378 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_385
timestamp 0
transform 1 0 20746 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_30_389
timestamp 0
transform 1 0 20930 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_30_391
timestamp 0
transform 1 0 21022 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_399
timestamp 0
transform 1 0 21390 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_407
timestamp 0
transform 1 0 21758 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_415
timestamp 0
transform 1 0 22126 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_423
timestamp 0
transform 1 0 22494 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_431
timestamp 0
transform 1 0 22862 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_439
timestamp 0
transform 1 0 23230 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_30_447
timestamp 0
transform 1 0 23598 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_30_449
timestamp 0
transform 1 0 23690 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_30_451
timestamp 0
transform 1 0 23782 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_459
timestamp 0
transform 1 0 24150 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_467
timestamp 0
transform 1 0 24518 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_475
timestamp 0
transform 1 0 24886 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_483
timestamp 0
transform 1 0 25254 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_491
timestamp 0
transform 1 0 25622 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_499
timestamp 0
transform 1 0 25990 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_30_507
timestamp 0
transform 1 0 26358 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_30_509
timestamp 0
transform 1 0 26450 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_30_511
timestamp 0
transform 1 0 26542 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_519
timestamp 0
transform 1 0 26910 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_527
timestamp 0
transform 1 0 27278 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_535
timestamp 0
transform 1 0 27646 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_543
timestamp 0
transform 1 0 28014 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_551
timestamp 0
transform 1 0 28382 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_30_559
timestamp 0
transform 1 0 28750 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_30_567
timestamp 0
transform 1 0 29118 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_30_569
timestamp 0
transform 1 0 29210 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_30_571
timestamp 0
transform 1 0 29302 0 1 11424
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_30_579
timestamp 0
transform 1 0 29670 0 1 11424
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_30_583
timestamp 0
transform 1 0 29854 0 1 11424
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_30_585
timestamp 0
transform 1 0 29946 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_31_0
timestamp 0
transform 1 0 3036 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_8
timestamp 0
transform 1 0 3404 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_16
timestamp 0
transform 1 0 3772 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_24
timestamp 0
transform 1 0 4140 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_32
timestamp 0
transform 1 0 4508 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_31_40
timestamp 0
transform 1 0 4876 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_31_44
timestamp 0
transform 1 0 5060 0 -1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_31_46
timestamp 0
transform 1 0 5152 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_31_56
timestamp 0
transform 1 0 5612 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_61
timestamp 0
transform 1 0 5842 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_31_65
timestamp 0
transform 1 0 6026 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_31_88
timestamp 0
transform 1 0 7084 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_116
timestamp 0
transform 1 0 8372 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_121
timestamp 0
transform 1 0 8602 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_31_125
timestamp 0
transform 1 0 8786 0 -1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_31_127
timestamp 0
transform 1 0 8878 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_31_135
timestamp 0
transform 1 0 9246 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_146
timestamp 0
transform 1 0 9752 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_174
timestamp 0
transform 1 0 11040 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_31_178
timestamp 0
transform 1 0 11224 0 -1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_31_181
timestamp 0
transform 1 0 11362 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 0
transform 1 0 11730 0 -1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_31_191
timestamp 0
transform 1 0 11822 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_31_208
timestamp 0
transform 1 0 12604 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_236
timestamp 0
transform 1 0 13892 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_241
timestamp 0
transform 1 0 14122 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_31_251
timestamp 0
transform 1 0 14582 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_259
timestamp 0
transform 1 0 14950 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_267
timestamp 0
transform 1 0 15318 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_275
timestamp 0
transform 1 0 15686 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_291
timestamp 0
transform 1 0 16422 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_31_299
timestamp 0
transform 1 0 16790 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_31_301
timestamp 0
transform 1 0 16882 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_309
timestamp 0
transform 1 0 17250 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_317
timestamp 0
transform 1 0 17618 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_325
timestamp 0
transform 1 0 17986 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_31_333
timestamp 0
transform 1 0 18354 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 0
transform 1 0 18538 0 -1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_31_339
timestamp 0
transform 1 0 18630 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_31_356
timestamp 0
transform 1 0 19412 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_31_361
timestamp 0
transform 1 0 19642 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_31_369
timestamp 0
transform 1 0 20010 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_31_397
timestamp 0
transform 1 0 21298 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_31_401
timestamp 0
transform 1 0 21482 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_31_408
timestamp 0
transform 1 0 21804 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_31_416
timestamp 0
transform 1 0 22172 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_31_421
timestamp 0
transform 1 0 22402 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_429
timestamp 0
transform 1 0 22770 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_437
timestamp 0
transform 1 0 23138 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_445
timestamp 0
transform 1 0 23506 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_453
timestamp 0
transform 1 0 23874 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_461
timestamp 0
transform 1 0 24242 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_469
timestamp 0
transform 1 0 24610 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_31_477
timestamp 0
transform 1 0 24978 0 -1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_31_479
timestamp 0
transform 1 0 25070 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_31_481
timestamp 0
transform 1 0 25162 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_489
timestamp 0
transform 1 0 25530 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_521
timestamp 0
transform 1 0 27002 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_529
timestamp 0
transform 1 0 27370 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_31_537
timestamp 0
transform 1 0 27738 0 -1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_31_539
timestamp 0
transform 1 0 27830 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_31_541
timestamp 0
transform 1 0 27922 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_549
timestamp 0
transform 1 0 28290 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_557
timestamp 0
transform 1 0 28658 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_565
timestamp 0
transform 1 0 29026 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_31_573
timestamp 0
transform 1 0 29394 0 -1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_31_581
timestamp 0
transform 1 0 29762 0 -1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_31_585
timestamp 0
transform 1 0 29946 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_32_0
timestamp 0
transform 1 0 3036 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_8
timestamp 0
transform 1 0 3404 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_16
timestamp 0
transform 1 0 3772 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_24
timestamp 0
transform 1 0 4140 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_28
timestamp 0
transform 1 0 4324 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_32_31
timestamp 0
transform 1 0 4462 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 0
transform 1 0 4646 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_56
timestamp 0
transform 1 0 5612 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_32_84
timestamp 0
transform 1 0 6900 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 0
transform 1 0 7084 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_32_91
timestamp 0
transform 1 0 7222 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_102
timestamp 0
transform 1 0 7728 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_110
timestamp 0
transform 1 0 8096 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_32_118
timestamp 0
transform 1 0 8464 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_143
timestamp 0
transform 1 0 9614 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_147
timestamp 0
transform 1 0 9798 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_149
timestamp 0
transform 1 0 9890 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_151
timestamp 0
transform 1 0 9982 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_179
timestamp 0
transform 1 0 11270 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_187
timestamp 0
transform 1 0 11638 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_197
timestamp 0
transform 1 0 12098 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_205
timestamp 0
transform 1 0 12466 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 0
transform 1 0 12650 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_211
timestamp 0
transform 1 0 12742 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_32_239
timestamp 0
transform 1 0 14030 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_32_249
timestamp 0
transform 1 0 14490 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 0
transform 1 0 14674 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_255
timestamp 0
transform 1 0 14766 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_32_259
timestamp 0
transform 1 0 14950 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_32_267
timestamp 0
transform 1 0 15318 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_269
timestamp 0
transform 1 0 15410 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_271
timestamp 0
transform 1 0 15502 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_275
timestamp 0
transform 1 0 15686 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_32_281
timestamp 0
transform 1 0 15962 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_288
timestamp 0
transform 1 0 16284 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_296
timestamp 0
transform 1 0 16652 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_300
timestamp 0
transform 1 0 16836 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_302
timestamp 0
transform 1 0 16928 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_306
timestamp 0
transform 1 0 17112 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_310
timestamp 0
transform 1 0 17296 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_32_317
timestamp 0
transform 1 0 17618 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_325
timestamp 0
transform 1 0 17986 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_32_329
timestamp 0
transform 1 0 18170 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_331
timestamp 0
transform 1 0 18262 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_342
timestamp 0
transform 1 0 18768 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_350
timestamp 0
transform 1 0 19136 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_354
timestamp 0
transform 1 0 19320 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_356
timestamp 0
transform 1 0 19412 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_361
timestamp 0
transform 1 0 19642 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_369
timestamp 0
transform 1 0 20010 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_377
timestamp 0
transform 1 0 20378 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_385
timestamp 0
transform 1 0 20746 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_32_389
timestamp 0
transform 1 0 20930 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_32_391
timestamp 0
transform 1 0 21022 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_399
timestamp 0
transform 1 0 21390 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_407
timestamp 0
transform 1 0 21758 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_415
timestamp 0
transform 1 0 22126 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_423
timestamp 0
transform 1 0 22494 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_431
timestamp 0
transform 1 0 22862 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_439
timestamp 0
transform 1 0 23230 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_32_447
timestamp 0
transform 1 0 23598 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_449
timestamp 0
transform 1 0 23690 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_32_451
timestamp 0
transform 1 0 23782 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_459
timestamp 0
transform 1 0 24150 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_467
timestamp 0
transform 1 0 24518 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_475
timestamp 0
transform 1 0 24886 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_479
timestamp 0
transform 1 0 25070 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_481
timestamp 0
transform 1 0 25162 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_32_506
timestamp 0
transform 1 0 26312 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_32_511
timestamp 0
transform 1 0 26542 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_519
timestamp 0
transform 1 0 26910 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_527
timestamp 0
transform 1 0 27278 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_535
timestamp 0
transform 1 0 27646 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_543
timestamp 0
transform 1 0 28014 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_551
timestamp 0
transform 1 0 28382 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_32_559
timestamp 0
transform 1 0 28750 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_32_567
timestamp 0
transform 1 0 29118 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_569
timestamp 0
transform 1 0 29210 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_32_571
timestamp 0
transform 1 0 29302 0 1 11968
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_32_579
timestamp 0
transform 1 0 29670 0 1 11968
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_32_583
timestamp 0
transform 1 0 29854 0 1 11968
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_32_585
timestamp 0
transform 1 0 29946 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_33_0
timestamp 0
transform 1 0 3036 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_8
timestamp 0
transform 1 0 3404 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_16
timestamp 0
transform 1 0 3772 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_24
timestamp 0
transform 1 0 4140 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_33_56
timestamp 0
transform 1 0 5612 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_33_61
timestamp 0
transform 1 0 5842 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_69
timestamp 0
transform 1 0 6210 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_33_77
timestamp 0
transform 1 0 6578 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_33_81
timestamp 0
transform 1 0 6762 0 -1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_33_107
timestamp 0
transform 1 0 7958 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_33_115
timestamp 0
transform 1 0 8326 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 0
transform 1 0 8510 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_33_121
timestamp 0
transform 1 0 8602 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_33_149
timestamp 0
transform 1 0 9890 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_33_175
timestamp 0
transform 1 0 11086 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_33_179
timestamp 0
transform 1 0 11270 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_33_181
timestamp 0
transform 1 0 11362 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_33_191
timestamp 0
transform 1 0 11822 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_33_200
timestamp 0
transform 1 0 12236 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 0
transform 1 0 12420 0 -1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_33_206
timestamp 0
transform 1 0 12512 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_33_231
timestamp 0
transform 1 0 13662 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_33_239
timestamp 0
transform 1 0 14030 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_33_241
timestamp 0
transform 1 0 14122 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_33_269
timestamp 0
transform 1 0 15410 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_33_289
timestamp 0
transform 1 0 16330 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 0
transform 1 0 16698 0 -1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_33_299
timestamp 0
transform 1 0 16790 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_33_301
timestamp 0
transform 1 0 16882 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_33_311
timestamp 0
transform 1 0 17342 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_33_319
timestamp 0
transform 1 0 17710 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_33_324
timestamp 0
transform 1 0 17940 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_336
timestamp 0
transform 1 0 18492 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_33_344
timestamp 0
transform 1 0 18860 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_33_348
timestamp 0
transform 1 0 19044 0 -1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_33_354
timestamp 0
transform 1 0 19320 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_33_358
timestamp 0
transform 1 0 19504 0 -1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_33_361
timestamp 0
transform 1 0 19642 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_369
timestamp 0
transform 1 0 20010 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_377
timestamp 0
transform 1 0 20378 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_385
timestamp 0
transform 1 0 20746 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_393
timestamp 0
transform 1 0 21114 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_401
timestamp 0
transform 1 0 21482 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_409
timestamp 0
transform 1 0 21850 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_33_417
timestamp 0
transform 1 0 22218 0 -1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_33_419
timestamp 0
transform 1 0 22310 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_33_421
timestamp 0
transform 1 0 22402 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_429
timestamp 0
transform 1 0 22770 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_437
timestamp 0
transform 1 0 23138 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_445
timestamp 0
transform 1 0 23506 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_458
timestamp 0
transform 1 0 24104 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_466
timestamp 0
transform 1 0 24472 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_33_474
timestamp 0
transform 1 0 24840 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_33_478
timestamp 0
transform 1 0 25024 0 -1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_33_481
timestamp 0
transform 1 0 25162 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_33_509
timestamp 0
transform 1 0 26450 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_33_520
timestamp 0
transform 1 0 26956 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_33_531
timestamp 0
transform 1 0 27462 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_33_539
timestamp 0
transform 1 0 27830 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_33_541
timestamp 0
transform 1 0 27922 0 -1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_33_569
timestamp 0
transform 1 0 29210 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_33_577
timestamp 0
transform 1 0 29578 0 -1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_33_585
timestamp 0
transform 1 0 29946 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_34_0
timestamp 0
transform 1 0 3036 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_34_26
timestamp 0
transform 1 0 4232 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_34_31
timestamp 0
transform 1 0 4462 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_39
timestamp 0
transform 1 0 4830 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_34_71
timestamp 0
transform 1 0 6302 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_34_79
timestamp 0
transform 1 0 6670 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_34_87
timestamp 0
transform 1 0 7038 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 0
transform 1 0 7130 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_91
timestamp 0
transform 1 0 7222 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_99
timestamp 0
transform 1 0 7590 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_34_107
timestamp 0
transform 1 0 7958 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_109
timestamp 0
transform 1 0 8050 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_134
timestamp 0
transform 1 0 9200 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_142
timestamp 0
transform 1 0 9568 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_151
timestamp 0
transform 1 0 9982 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_159
timestamp 0
transform 1 0 10350 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_34_167
timestamp 0
transform 1 0 10718 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 0
transform 1 0 10810 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_194
timestamp 0
transform 1 0 11960 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_202
timestamp 0
transform 1 0 12328 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_211
timestamp 0
transform 1 0 12742 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_219
timestamp 0
transform 1 0 13110 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_227
timestamp 0
transform 1 0 13478 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_34_235
timestamp 0
transform 1 0 13846 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_241
timestamp 0
transform 1 0 14122 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_254
timestamp 0
transform 1 0 14720 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_262
timestamp 0
transform 1 0 15088 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_34_271
timestamp 0
transform 1 0 15502 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_34_278
timestamp 0
transform 1 0 15824 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_34_286
timestamp 0
transform 1 0 16192 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_34_299
timestamp 0
transform 1 0 16790 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_307
timestamp 0
transform 1 0 17158 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_315
timestamp 0
transform 1 0 17526 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_34_323
timestamp 0
transform 1 0 17894 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_34_327
timestamp 0
transform 1 0 18078 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_329
timestamp 0
transform 1 0 18170 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_331
timestamp 0
transform 1 0 18262 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_339
timestamp 0
transform 1 0 18630 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_347
timestamp 0
transform 1 0 18998 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_355
timestamp 0
transform 1 0 19366 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_34_363
timestamp 0
transform 1 0 19734 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_34_367
timestamp 0
transform 1 0 19918 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 0
transform 1 0 20010 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_379
timestamp 0
transform 1 0 20470 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_34_387
timestamp 0
transform 1 0 20838 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_389
timestamp 0
transform 1 0 20930 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_34_391
timestamp 0
transform 1 0 21022 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_34_419
timestamp 0
transform 1 0 22310 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_427
timestamp 0
transform 1 0 22678 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_435
timestamp 0
transform 1 0 23046 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_34_443
timestamp 0
transform 1 0 23414 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_34_447
timestamp 0
transform 1 0 23598 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_449
timestamp 0
transform 1 0 23690 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_451
timestamp 0
transform 1 0 23782 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_459
timestamp 0
transform 1 0 24150 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_467
timestamp 0
transform 1 0 24518 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_475
timestamp 0
transform 1 0 24886 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_483
timestamp 0
transform 1 0 25254 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_491
timestamp 0
transform 1 0 25622 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_499
timestamp 0
transform 1 0 25990 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_34_507
timestamp 0
transform 1 0 26358 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_509
timestamp 0
transform 1 0 26450 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_511
timestamp 0
transform 1 0 26542 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_519
timestamp 0
transform 1 0 26910 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_34_527
timestamp 0
transform 1 0 27278 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_34_535
timestamp 0
transform 1 0 27646 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_34_563
timestamp 0
transform 1 0 28934 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_34_567
timestamp 0
transform 1 0 29118 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_569
timestamp 0
transform 1 0 29210 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_34_571
timestamp 0
transform 1 0 29302 0 1 12512
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_34_579
timestamp 0
transform 1 0 29670 0 1 12512
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_34_583
timestamp 0
transform 1 0 29854 0 1 12512
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_34_585
timestamp 0
transform 1 0 29946 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_35_0
timestamp 0
transform 1 0 3036 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_8
timestamp 0
transform 1 0 3404 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_35_12
timestamp 0
transform 1 0 3588 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_35_37
timestamp 0
transform 1 0 4738 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_45
timestamp 0
transform 1 0 5106 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_53
timestamp 0
transform 1 0 5474 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 0
transform 1 0 5658 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_35_59
timestamp 0
transform 1 0 5750 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_35_61
timestamp 0
transform 1 0 5842 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 0
transform 1 0 6026 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_35_67
timestamp 0
transform 1 0 6118 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_35_75
timestamp 0
transform 1 0 6486 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_35_83
timestamp 0
transform 1 0 6854 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_35_109
timestamp 0
transform 1 0 8050 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_35_117
timestamp 0
transform 1 0 8418 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 0
transform 1 0 8510 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_35_121
timestamp 0
transform 1 0 8602 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_129
timestamp 0
transform 1 0 8970 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_137
timestamp 0
transform 1 0 9338 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_145
timestamp 0
transform 1 0 9706 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 0
transform 1 0 9890 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_35_151
timestamp 0
transform 1 0 9982 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_35_176
timestamp 0
transform 1 0 11132 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_35_181
timestamp 0
transform 1 0 11362 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_197
timestamp 0
transform 1 0 12098 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_35_206
timestamp 0
transform 1 0 12512 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 0
transform 1 0 12696 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_35_236
timestamp 0
transform 1 0 13892 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_35_241
timestamp 0
transform 1 0 14122 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_249
timestamp 0
transform 1 0 14490 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_257
timestamp 0
transform 1 0 14858 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_265
timestamp 0
transform 1 0 15226 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_273
timestamp 0
transform 1 0 15594 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_281
timestamp 0
transform 1 0 15962 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_35_296
timestamp 0
transform 1 0 16652 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_35_301
timestamp 0
transform 1 0 16882 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_309
timestamp 0
transform 1 0 17250 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_317
timestamp 0
transform 1 0 17618 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_325
timestamp 0
transform 1 0 17986 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_333
timestamp 0
transform 1 0 18354 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_341
timestamp 0
transform 1 0 18722 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_35_349
timestamp 0
transform 1 0 19090 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_35_356
timestamp 0
transform 1 0 19412 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_35_361
timestamp 0
transform 1 0 19642 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_369
timestamp 0
transform 1 0 20010 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_377
timestamp 0
transform 1 0 20378 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_35_385
timestamp 0
transform 1 0 20746 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_35_410
timestamp 0
transform 1 0 21896 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_35_418
timestamp 0
transform 1 0 22264 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_35_421
timestamp 0
transform 1 0 22402 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_35_433
timestamp 0
transform 1 0 22954 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_441
timestamp 0
transform 1 0 23322 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_449
timestamp 0
transform 1 0 23690 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_457
timestamp 0
transform 1 0 24058 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_465
timestamp 0
transform 1 0 24426 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_473
timestamp 0
transform 1 0 24794 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_477
timestamp 0
transform 1 0 24978 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_35_479
timestamp 0
transform 1 0 25070 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_35_481
timestamp 0
transform 1 0 25162 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_489
timestamp 0
transform 1 0 25530 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_493
timestamp 0
transform 1 0 25714 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_35_495
timestamp 0
transform 1 0 25806 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_35_520
timestamp 0
transform 1 0 26956 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_35_528
timestamp 0
transform 1 0 27324 0 -1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_35_536
timestamp 0
transform 1 0 27692 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_35_541
timestamp 0
transform 1 0 27922 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_545
timestamp 0
transform 1 0 28106 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_35_571
timestamp 0
transform 1 0 29302 0 -1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_35_583
timestamp 0
transform 1 0 29854 0 -1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_35_585
timestamp 0
transform 1 0 29946 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_36_0
timestamp 0
transform 1 0 3036 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_36_26
timestamp 0
transform 1 0 4232 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_36_31
timestamp 0
transform 1 0 4462 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_36_41
timestamp 0
transform 1 0 4922 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_36_49
timestamp 0
transform 1 0 5290 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_36_74
timestamp 0
transform 1 0 6440 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_82
timestamp 0
transform 1 0 6808 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_91
timestamp 0
transform 1 0 7222 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_36_99
timestamp 0
transform 1 0 7590 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_36_103
timestamp 0
transform 1 0 7774 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_36_113
timestamp 0
transform 1 0 8234 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_36_121
timestamp 0
transform 1 0 8602 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_36_146
timestamp 0
transform 1 0 9752 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_36_151
timestamp 0
transform 1 0 9982 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_159
timestamp 0
transform 1 0 10350 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_167
timestamp 0
transform 1 0 10718 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_36_175
timestamp 0
transform 1 0 11086 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_36_179
timestamp 0
transform 1 0 11270 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_36_181
timestamp 0
transform 1 0 11362 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_36_206
timestamp 0
transform 1 0 12512 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_36_211
timestamp 0
transform 1 0 12742 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 0
transform 1 0 13110 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_36_221
timestamp 0
transform 1 0 13202 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_36_246
timestamp 0
transform 1 0 14352 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_36_258
timestamp 0
transform 1 0 14904 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_36_266
timestamp 0
transform 1 0 15272 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_36_271
timestamp 0
transform 1 0 15502 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_36_279
timestamp 0
transform 1 0 15870 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_36_285
timestamp 0
transform 1 0 16146 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_36_293
timestamp 0
transform 1 0 16514 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_301
timestamp 0
transform 1 0 16882 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_309
timestamp 0
transform 1 0 17250 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_317
timestamp 0
transform 1 0 17618 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_36_325
timestamp 0
transform 1 0 17986 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_36_329
timestamp 0
transform 1 0 18170 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_36_331
timestamp 0
transform 1 0 18262 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_343
timestamp 0
transform 1 0 18814 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_351
timestamp 0
transform 1 0 19182 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_359
timestamp 0
transform 1 0 19550 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_367
timestamp 0
transform 1 0 19918 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_375
timestamp 0
transform 1 0 20286 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_36_383
timestamp 0
transform 1 0 20654 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_36_387
timestamp 0
transform 1 0 20838 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_36_389
timestamp 0
transform 1 0 20930 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_36_391
timestamp 0
transform 1 0 21022 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_36_419
timestamp 0
transform 1 0 22310 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_427
timestamp 0
transform 1 0 22678 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_435
timestamp 0
transform 1 0 23046 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_36_443
timestamp 0
transform 1 0 23414 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_36_447
timestamp 0
transform 1 0 23598 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_36_449
timestamp 0
transform 1 0 23690 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_36_451
timestamp 0
transform 1 0 23782 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_459
timestamp 0
transform 1 0 24150 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_467
timestamp 0
transform 1 0 24518 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_475
timestamp 0
transform 1 0 24886 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_483
timestamp 0
transform 1 0 25254 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_491
timestamp 0
transform 1 0 25622 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_499
timestamp 0
transform 1 0 25990 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_36_507
timestamp 0
transform 1 0 26358 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_36_509
timestamp 0
transform 1 0 26450 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_36_511
timestamp 0
transform 1 0 26542 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_519
timestamp 0
transform 1 0 26910 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_527
timestamp 0
transform 1 0 27278 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_535
timestamp 0
transform 1 0 27646 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_543
timestamp 0
transform 1 0 28014 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_551
timestamp 0
transform 1 0 28382 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_36_559
timestamp 0
transform 1 0 28750 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_36_567
timestamp 0
transform 1 0 29118 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_36_569
timestamp 0
transform 1 0 29210 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_36_571
timestamp 0
transform 1 0 29302 0 1 13056
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_36_579
timestamp 0
transform 1 0 29670 0 1 13056
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_36_583
timestamp 0
transform 1 0 29854 0 1 13056
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_36_585
timestamp 0
transform 1 0 29946 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_37_0
timestamp 0
transform 1 0 3036 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_37_4
timestamp 0
transform 1 0 3220 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_37_30
timestamp 0
transform 1 0 4416 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_37_40
timestamp 0
transform 1 0 4876 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_37_48
timestamp 0
transform 1 0 5244 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_37_56
timestamp 0
transform 1 0 5612 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_37_61
timestamp 0
transform 1 0 5842 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_69
timestamp 0
transform 1 0 6210 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_37_77
timestamp 0
transform 1 0 6578 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_37_81
timestamp 0
transform 1 0 6762 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_37_83
timestamp 0
transform 1 0 6854 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_37_108
timestamp 0
transform 1 0 8004 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_37_116
timestamp 0
transform 1 0 8372 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_37_121
timestamp 0
transform 1 0 8602 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_37_129
timestamp 0
transform 1 0 8970 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_37_136
timestamp 0
transform 1 0 9292 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_37_147
timestamp 0
transform 1 0 9798 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_37_151
timestamp 0
transform 1 0 9982 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_37_176
timestamp 0
transform 1 0 11132 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_37_181
timestamp 0
transform 1 0 11362 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_189
timestamp 0
transform 1 0 11730 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_37_197
timestamp 0
transform 1 0 12098 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_37_201
timestamp 0
transform 1 0 12282 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_37_205
timestamp 0
transform 1 0 12466 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_37_209
timestamp 0
transform 1 0 12650 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_37_211
timestamp 0
transform 1 0 12742 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_37_236
timestamp 0
transform 1 0 13892 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_37_241
timestamp 0
transform 1 0 14122 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_37_269
timestamp 0
transform 1 0 15410 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_37_289
timestamp 0
transform 1 0 16330 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_37_297
timestamp 0
transform 1 0 16698 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_37_299
timestamp 0
transform 1 0 16790 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_37_301
timestamp 0
transform 1 0 16882 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_309
timestamp 0
transform 1 0 17250 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_317
timestamp 0
transform 1 0 17618 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_325
timestamp 0
transform 1 0 17986 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_37_333
timestamp 0
transform 1 0 18354 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_37_339
timestamp 0
transform 1 0 18630 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_37_349
timestamp 0
transform 1 0 19090 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_37_357
timestamp 0
transform 1 0 19458 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_37_359
timestamp 0
transform 1 0 19550 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_37_361
timestamp 0
transform 1 0 19642 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_369
timestamp 0
transform 1 0 20010 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_377
timestamp 0
transform 1 0 20378 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_385
timestamp 0
transform 1 0 20746 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_393
timestamp 0
transform 1 0 21114 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_401
timestamp 0
transform 1 0 21482 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_409
timestamp 0
transform 1 0 21850 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_37_417
timestamp 0
transform 1 0 22218 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_37_419
timestamp 0
transform 1 0 22310 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_37_421
timestamp 0
transform 1 0 22402 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_429
timestamp 0
transform 1 0 22770 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_437
timestamp 0
transform 1 0 23138 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_445
timestamp 0
transform 1 0 23506 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_37_453
timestamp 0
transform 1 0 23874 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_37_457
timestamp 0
transform 1 0 24058 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_37_463
timestamp 0
transform 1 0 24334 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_471
timestamp 0
transform 1 0 24702 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_37_479
timestamp 0
transform 1 0 25070 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_37_481
timestamp 0
transform 1 0 25162 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_489
timestamp 0
transform 1 0 25530 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_37_497
timestamp 0
transform 1 0 25898 0 -1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_37_523
timestamp 0
transform 1 0 27094 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_531
timestamp 0
transform 1 0 27462 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_37_539
timestamp 0
transform 1 0 27830 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_37_541
timestamp 0
transform 1 0 27922 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_549
timestamp 0
transform 1 0 28290 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_557
timestamp 0
transform 1 0 28658 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_565
timestamp 0
transform 1 0 29026 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_37_573
timestamp 0
transform 1 0 29394 0 -1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_37_581
timestamp 0
transform 1 0 29762 0 -1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_37_585
timestamp 0
transform 1 0 29946 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_0
timestamp 0
transform 1 0 3036 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_8
timestamp 0
transform 1 0 3404 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_16
timestamp 0
transform 1 0 3772 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_24
timestamp 0
transform 1 0 4140 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_38_28
timestamp 0
transform 1 0 4324 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_38_31
timestamp 0
transform 1 0 4462 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_39
timestamp 0
transform 1 0 4830 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_38_43
timestamp 0
transform 1 0 5014 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 0
transform 1 0 5106 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_70
timestamp 0
transform 1 0 6256 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_78
timestamp 0
transform 1 0 6624 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_86
timestamp 0
transform 1 0 6992 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_38_91
timestamp 0
transform 1 0 7222 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_99
timestamp 0
transform 1 0 7590 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_107
timestamp 0
transform 1 0 7958 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_38_115
timestamp 0
transform 1 0 8326 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_38_117
timestamp 0
transform 1 0 8418 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_142
timestamp 0
transform 1 0 9568 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_151
timestamp 0
transform 1 0 9982 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_159
timestamp 0
transform 1 0 10350 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_38_163
timestamp 0
transform 1 0 10534 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_38_165
timestamp 0
transform 1 0 10626 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_190
timestamp 0
transform 1 0 11776 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_198
timestamp 0
transform 1 0 12144 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_206
timestamp 0
transform 1 0 12512 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_38_211
timestamp 0
transform 1 0 12742 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_219
timestamp 0
transform 1 0 13110 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_227
timestamp 0
transform 1 0 13478 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_235
timestamp 0
transform 1 0 13846 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_38_239
timestamp 0
transform 1 0 14030 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_38_241
timestamp 0
transform 1 0 14122 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_38_266
timestamp 0
transform 1 0 15272 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_38_271
timestamp 0
transform 1 0 15502 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_279
timestamp 0
transform 1 0 15870 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_287
timestamp 0
transform 1 0 16238 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_38_295
timestamp 0
transform 1 0 16606 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_300
timestamp 0
transform 1 0 16836 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_308
timestamp 0
transform 1 0 17204 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_316
timestamp 0
transform 1 0 17572 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_324
timestamp 0
transform 1 0 17940 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_38_328
timestamp 0
transform 1 0 18124 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_38_331
timestamp 0
transform 1 0 18262 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_38_339
timestamp 0
transform 1 0 18630 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_356
timestamp 0
transform 1 0 19412 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_364
timestamp 0
transform 1 0 19780 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_372
timestamp 0
transform 1 0 20148 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_380
timestamp 0
transform 1 0 20516 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_38_388
timestamp 0
transform 1 0 20884 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_38_391
timestamp 0
transform 1 0 21022 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_399
timestamp 0
transform 1 0 21390 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_407
timestamp 0
transform 1 0 21758 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_415
timestamp 0
transform 1 0 22126 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_423
timestamp 0
transform 1 0 22494 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_38_431
timestamp 0
transform 1 0 22862 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_38_433
timestamp 0
transform 1 0 22954 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_438
timestamp 0
transform 1 0 23184 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_446
timestamp 0
transform 1 0 23552 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_38_451
timestamp 0
transform 1 0 23782 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_459
timestamp 0
transform 1 0 24150 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_38_463
timestamp 0
transform 1 0 24334 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_38_465
timestamp 0
transform 1 0 24426 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_490
timestamp 0
transform 1 0 25576 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_498
timestamp 0
transform 1 0 25944 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_506
timestamp 0
transform 1 0 26312 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_38_511
timestamp 0
transform 1 0 26542 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_38_515
timestamp 0
transform 1 0 26726 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_521
timestamp 0
transform 1 0 27002 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_529
timestamp 0
transform 1 0 27370 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_537
timestamp 0
transform 1 0 27738 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_38_545
timestamp 0
transform 1 0 28106 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_38_553
timestamp 0
transform 1 0 28474 0 1 13600
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_38_555
timestamp 0
transform 1 0 28566 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_38_562
timestamp 0
transform 1 0 28888 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_38_571
timestamp 0
transform 1 0 29302 0 1 13600
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_38_578
timestamp 0
transform 1 0 29624 0 1 13600
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_0
timestamp 0
transform 1 0 3036 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_8
timestamp 0
transform 1 0 3404 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_16
timestamp 0
transform 1 0 3772 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_24
timestamp 0
transform 1 0 4140 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_39_56
timestamp 0
transform 1 0 5612 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_39_61
timestamp 0
transform 1 0 5842 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_39_65
timestamp 0
transform 1 0 6026 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_39_74
timestamp 0
transform 1 0 6440 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_82
timestamp 0
transform 1 0 6808 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_90
timestamp 0
transform 1 0 7176 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_98
timestamp 0
transform 1 0 7544 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_106
timestamp 0
transform 1 0 7912 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_39_114
timestamp 0
transform 1 0 8280 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 0
transform 1 0 8464 0 -1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_39_121
timestamp 0
transform 1 0 8602 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_129
timestamp 0
transform 1 0 8970 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_39_137
timestamp 0
transform 1 0 9338 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_39_141
timestamp 0
transform 1 0 9522 0 -1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_39_149
timestamp 0
transform 1 0 9890 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_157
timestamp 0
transform 1 0 10258 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_165
timestamp 0
transform 1 0 10626 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_39_173
timestamp 0
transform 1 0 10994 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_39_177
timestamp 0
transform 1 0 11178 0 -1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_39_179
timestamp 0
transform 1 0 11270 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_39_181
timestamp 0
transform 1 0 11362 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_189
timestamp 0
transform 1 0 11730 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_197
timestamp 0
transform 1 0 12098 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_205
timestamp 0
transform 1 0 12466 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_213
timestamp 0
transform 1 0 12834 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_221
timestamp 0
transform 1 0 13202 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_229
timestamp 0
transform 1 0 13570 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_39_237
timestamp 0
transform 1 0 13938 0 -1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_39_239
timestamp 0
transform 1 0 14030 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_39_241
timestamp 0
transform 1 0 14122 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_249
timestamp 0
transform 1 0 14490 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_257
timestamp 0
transform 1 0 14858 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_272
timestamp 0
transform 1 0 15548 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_280
timestamp 0
transform 1 0 15916 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_288
timestamp 0
transform 1 0 16284 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_39_296
timestamp 0
transform 1 0 16652 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_39_301
timestamp 0
transform 1 0 16882 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_39_321
timestamp 0
transform 1 0 17802 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_329
timestamp 0
transform 1 0 18170 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_337
timestamp 0
transform 1 0 18538 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_345
timestamp 0
transform 1 0 18906 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_39_353
timestamp 0
transform 1 0 19274 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_39_357
timestamp 0
transform 1 0 19458 0 -1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_39_359
timestamp 0
transform 1 0 19550 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_39_361
timestamp 0
transform 1 0 19642 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_39_376
timestamp 0
transform 1 0 20332 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_39_385
timestamp 0
transform 1 0 20746 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_39_393
timestamp 0
transform 1 0 21114 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_39_397
timestamp 0
transform 1 0 21298 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_39_403
timestamp 0
transform 1 0 21574 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_411
timestamp 0
transform 1 0 21942 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_39_419
timestamp 0
transform 1 0 22310 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_39_421
timestamp 0
transform 1 0 22402 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_429
timestamp 0
transform 1 0 22770 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_437
timestamp 0
transform 1 0 23138 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_445
timestamp 0
transform 1 0 23506 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_453
timestamp 0
transform 1 0 23874 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_461
timestamp 0
transform 1 0 24242 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_469
timestamp 0
transform 1 0 24610 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_39_477
timestamp 0
transform 1 0 24978 0 -1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_39_479
timestamp 0
transform 1 0 25070 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_39_481
timestamp 0
transform 1 0 25162 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_489
timestamp 0
transform 1 0 25530 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_39_497
timestamp 0
transform 1 0 25898 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_39_522
timestamp 0
transform 1 0 27048 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_39_534
timestamp 0
transform 1 0 27600 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_39_538
timestamp 0
transform 1 0 27784 0 -1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_39_541
timestamp 0
transform 1 0 27922 0 -1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_39_569
timestamp 0
transform 1 0 29210 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_39_577
timestamp 0
transform 1 0 29578 0 -1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_39_585
timestamp 0
transform 1 0 29946 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_40_0
timestamp 0
transform 1 0 3036 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_40_26
timestamp 0
transform 1 0 4232 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_40_31
timestamp 0
transform 1 0 4462 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_39
timestamp 0
transform 1 0 4830 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_47
timestamp 0
transform 1 0 5198 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_40_55
timestamp 0
transform 1 0 5566 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_40_83
timestamp 0
transform 1 0 6854 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_40_87
timestamp 0
transform 1 0 7038 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 0
transform 1 0 7130 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_91
timestamp 0
transform 1 0 7222 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_40_99
timestamp 0
transform 1 0 7590 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_124
timestamp 0
transform 1 0 8740 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_132
timestamp 0
transform 1 0 9108 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_140
timestamp 0
transform 1 0 9476 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_40_148
timestamp 0
transform 1 0 9844 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_40_151
timestamp 0
transform 1 0 9982 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_159
timestamp 0
transform 1 0 10350 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_40_167
timestamp 0
transform 1 0 10718 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_169
timestamp 0
transform 1 0 10810 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_40_194
timestamp 0
transform 1 0 11960 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_40_205
timestamp 0
transform 1 0 12466 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_40_209
timestamp 0
transform 1 0 12650 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_211
timestamp 0
transform 1 0 12742 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_40_219
timestamp 0
transform 1 0 13110 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_221
timestamp 0
transform 1 0 13202 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_246
timestamp 0
transform 1 0 14352 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_254
timestamp 0
transform 1 0 14720 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_262
timestamp 0
transform 1 0 15088 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_271
timestamp 0
transform 1 0 15502 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_279
timestamp 0
transform 1 0 15870 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_287
timestamp 0
transform 1 0 16238 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_295
timestamp 0
transform 1 0 16606 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_40_303
timestamp 0
transform 1 0 16974 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_40_307
timestamp 0
transform 1 0 17158 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_309
timestamp 0
transform 1 0 17250 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_40_314
timestamp 0
transform 1 0 17480 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_40_323
timestamp 0
transform 1 0 17894 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_40_327
timestamp 0
transform 1 0 18078 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_329
timestamp 0
transform 1 0 18170 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_331
timestamp 0
transform 1 0 18262 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_339
timestamp 0
transform 1 0 18630 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_347
timestamp 0
transform 1 0 18998 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_40_355
timestamp 0
transform 1 0 19366 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_40_368
timestamp 0
transform 1 0 19964 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_376
timestamp 0
transform 1 0 20332 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_40_384
timestamp 0
transform 1 0 20700 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_40_388
timestamp 0
transform 1 0 20884 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_40_391
timestamp 0
transform 1 0 21022 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_40_399
timestamp 0
transform 1 0 21390 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_407
timestamp 0
transform 1 0 21758 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_415
timestamp 0
transform 1 0 22126 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_423
timestamp 0
transform 1 0 22494 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_435
timestamp 0
transform 1 0 23046 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_40_443
timestamp 0
transform 1 0 23414 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_40_447
timestamp 0
transform 1 0 23598 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_449
timestamp 0
transform 1 0 23690 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_451
timestamp 0
transform 1 0 23782 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_40_459
timestamp 0
transform 1 0 24150 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_40_487
timestamp 0
transform 1 0 25438 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_40_499
timestamp 0
transform 1 0 25990 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_40_507
timestamp 0
transform 1 0 26358 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_509
timestamp 0
transform 1 0 26450 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_511
timestamp 0
transform 1 0 26542 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_519
timestamp 0
transform 1 0 26910 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_40_527
timestamp 0
transform 1 0 27278 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_40_535
timestamp 0
transform 1 0 27646 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_40_560
timestamp 0
transform 1 0 28796 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_40_568
timestamp 0
transform 1 0 29164 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_40_571
timestamp 0
transform 1 0 29302 0 1 14144
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_40_579
timestamp 0
transform 1 0 29670 0 1 14144
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_40_583
timestamp 0
transform 1 0 29854 0 1 14144
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_40_585
timestamp 0
transform 1 0 29946 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_0
timestamp 0
transform 1 0 3036 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_8
timestamp 0
transform 1 0 3404 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_40
timestamp 0
transform 1 0 4876 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_48
timestamp 0
transform 1 0 5244 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_56
timestamp 0
transform 1 0 5612 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_41_61
timestamp 0
transform 1 0 5842 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_69
timestamp 0
transform 1 0 6210 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 0
transform 1 0 6578 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_41_103
timestamp 0
transform 1 0 7774 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_111
timestamp 0
transform 1 0 8142 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_41_119
timestamp 0
transform 1 0 8510 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_121
timestamp 0
transform 1 0 8602 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_41_129
timestamp 0
transform 1 0 8970 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 0
transform 1 0 9062 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_156
timestamp 0
transform 1 0 10212 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_164
timestamp 0
transform 1 0 10580 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_172
timestamp 0
transform 1 0 10948 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_181
timestamp 0
transform 1 0 11362 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_189
timestamp 0
transform 1 0 11730 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_197
timestamp 0
transform 1 0 12098 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_41_201
timestamp 0
transform 1 0 12282 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_41_227
timestamp 0
transform 1 0 13478 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_235
timestamp 0
transform 1 0 13846 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_41_239
timestamp 0
transform 1 0 14030 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_241
timestamp 0
transform 1 0 14122 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_249
timestamp 0
transform 1 0 14490 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_257
timestamp 0
transform 1 0 14858 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_41_261
timestamp 0
transform 1 0 15042 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_41_263
timestamp 0
transform 1 0 15134 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_288
timestamp 0
transform 1 0 16284 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_296
timestamp 0
transform 1 0 16652 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_41_301
timestamp 0
transform 1 0 16882 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_309
timestamp 0
transform 1 0 17250 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_317
timestamp 0
transform 1 0 17618 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_325
timestamp 0
transform 1 0 17986 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_333
timestamp 0
transform 1 0 18354 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_341
timestamp 0
transform 1 0 18722 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_349
timestamp 0
transform 1 0 19090 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_41_357
timestamp 0
transform 1 0 19458 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_41_359
timestamp 0
transform 1 0 19550 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_361
timestamp 0
transform 1 0 19642 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_369
timestamp 0
transform 1 0 20010 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_377
timestamp 0
transform 1 0 20378 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_385
timestamp 0
transform 1 0 20746 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_393
timestamp 0
transform 1 0 21114 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_401
timestamp 0
transform 1 0 21482 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_409
timestamp 0
transform 1 0 21850 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_41_417
timestamp 0
transform 1 0 22218 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_41_419
timestamp 0
transform 1 0 22310 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_421
timestamp 0
transform 1 0 22402 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_429
timestamp 0
transform 1 0 22770 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_437
timestamp 0
transform 1 0 23138 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_445
timestamp 0
transform 1 0 23506 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_453
timestamp 0
transform 1 0 23874 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_461
timestamp 0
transform 1 0 24242 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_469
timestamp 0
transform 1 0 24610 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_41_477
timestamp 0
transform 1 0 24978 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_41_479
timestamp 0
transform 1 0 25070 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_481
timestamp 0
transform 1 0 25162 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_489
timestamp 0
transform 1 0 25530 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_497
timestamp 0
transform 1 0 25898 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_41_501
timestamp 0
transform 1 0 26082 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_41_527
timestamp 0
transform 1 0 27278 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_535
timestamp 0
transform 1 0 27646 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_41_539
timestamp 0
transform 1 0 27830 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_541
timestamp 0
transform 1 0 27922 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_549
timestamp 0
transform 1 0 28290 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_41_557
timestamp 0
transform 1 0 28658 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_41_565
timestamp 0
transform 1 0 29026 0 -1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_41_569
timestamp 0
transform 1 0 29210 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_41_571
timestamp 0
transform 1 0 29302 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_41_575
timestamp 0
transform 1 0 29486 0 -1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_41_583
timestamp 0
transform 1 0 29854 0 -1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_41_585
timestamp 0
transform 1 0 29946 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_42_0
timestamp 0
transform 1 0 3036 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_42_26
timestamp 0
transform 1 0 4232 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_42_31
timestamp 0
transform 1 0 4462 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_42_35
timestamp 0
transform 1 0 4646 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_42_44
timestamp 0
transform 1 0 5060 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_52
timestamp 0
transform 1 0 5428 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 0
transform 1 0 5796 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_42_86
timestamp 0
transform 1 0 6992 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_42_91
timestamp 0
transform 1 0 7222 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_42_102
timestamp 0
transform 1 0 7728 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_110
timestamp 0
transform 1 0 8096 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_42_118
timestamp 0
transform 1 0 8464 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_42_146
timestamp 0
transform 1 0 9752 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_42_151
timestamp 0
transform 1 0 9982 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_42_163
timestamp 0
transform 1 0 10534 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_171
timestamp 0
transform 1 0 10902 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_42_179
timestamp 0
transform 1 0 11270 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_42_181
timestamp 0
transform 1 0 11362 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_42_206
timestamp 0
transform 1 0 12512 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_42_211
timestamp 0
transform 1 0 12742 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_42_219
timestamp 0
transform 1 0 13110 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_42_223
timestamp 0
transform 1 0 13294 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_42_233
timestamp 0
transform 1 0 13754 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_42_241
timestamp 0
transform 1 0 14122 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_42_266
timestamp 0
transform 1 0 15272 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_42_271
timestamp 0
transform 1 0 15502 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_42_279
timestamp 0
transform 1 0 15870 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_42_286
timestamp 0
transform 1 0 16192 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_294
timestamp 0
transform 1 0 16560 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_302
timestamp 0
transform 1 0 16928 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_310
timestamp 0
transform 1 0 17296 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_318
timestamp 0
transform 1 0 17664 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_42_326
timestamp 0
transform 1 0 18032 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_42_331
timestamp 0
transform 1 0 18262 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_339
timestamp 0
transform 1 0 18630 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_347
timestamp 0
transform 1 0 18998 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_355
timestamp 0
transform 1 0 19366 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_363
timestamp 0
transform 1 0 19734 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_371
timestamp 0
transform 1 0 20102 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_379
timestamp 0
transform 1 0 20470 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_42_387
timestamp 0
transform 1 0 20838 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_42_389
timestamp 0
transform 1 0 20930 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_42_391
timestamp 0
transform 1 0 21022 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_399
timestamp 0
transform 1 0 21390 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_407
timestamp 0
transform 1 0 21758 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_415
timestamp 0
transform 1 0 22126 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_423
timestamp 0
transform 1 0 22494 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_431
timestamp 0
transform 1 0 22862 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_439
timestamp 0
transform 1 0 23230 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_42_447
timestamp 0
transform 1 0 23598 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_42_449
timestamp 0
transform 1 0 23690 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_42_451
timestamp 0
transform 1 0 23782 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_459
timestamp 0
transform 1 0 24150 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_42_467
timestamp 0
transform 1 0 24518 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_42_493
timestamp 0
transform 1 0 25714 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_501
timestamp 0
transform 1 0 26082 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_42_509
timestamp 0
transform 1 0 26450 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_42_511
timestamp 0
transform 1 0 26542 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_519
timestamp 0
transform 1 0 26910 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_527
timestamp 0
transform 1 0 27278 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_535
timestamp 0
transform 1 0 27646 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_543
timestamp 0
transform 1 0 28014 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_551
timestamp 0
transform 1 0 28382 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_42_559
timestamp 0
transform 1 0 28750 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_42_567
timestamp 0
transform 1 0 29118 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_42_569
timestamp 0
transform 1 0 29210 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_42_571
timestamp 0
transform 1 0 29302 0 1 14688
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_42_579
timestamp 0
transform 1 0 29670 0 1 14688
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_42_583
timestamp 0
transform 1 0 29854 0 1 14688
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_42_585
timestamp 0
transform 1 0 29946 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_43_0
timestamp 0
transform 1 0 3036 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_43_8
timestamp 0
transform 1 0 3404 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_10
timestamp 0
transform 1 0 3496 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_43_35
timestamp 0
transform 1 0 4646 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_43_46
timestamp 0
transform 1 0 5152 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_43_54
timestamp 0
transform 1 0 5520 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_43_58
timestamp 0
transform 1 0 5704 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_43_61
timestamp 0
transform 1 0 5842 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 0
transform 1 0 6210 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_71
timestamp 0
transform 1 0 6302 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_43_77
timestamp 0
transform 1 0 6578 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_43_88
timestamp 0
transform 1 0 7084 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_43_116
timestamp 0
transform 1 0 8372 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_43_121
timestamp 0
transform 1 0 8602 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_43_133
timestamp 0
transform 1 0 9154 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_141
timestamp 0
transform 1 0 9522 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_43_149
timestamp 0
transform 1 0 9890 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_151
timestamp 0
transform 1 0 9982 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_43_176
timestamp 0
transform 1 0 11132 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_43_181
timestamp 0
transform 1 0 11362 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_43_185
timestamp 0
transform 1 0 11546 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_187
timestamp 0
transform 1 0 11638 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_43_196
timestamp 0
transform 1 0 12052 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_204
timestamp 0
transform 1 0 12420 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_43_236
timestamp 0
transform 1 0 13892 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_43_241
timestamp 0
transform 1 0 14122 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_43_245
timestamp 0
transform 1 0 14306 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_247
timestamp 0
transform 1 0 14398 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_43_256
timestamp 0
transform 1 0 14812 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_43_264
timestamp 0
transform 1 0 15180 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_43_292
timestamp 0
transform 1 0 16468 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_301
timestamp 0
transform 1 0 16882 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_309
timestamp 0
transform 1 0 17250 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_317
timestamp 0
transform 1 0 17618 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_325
timestamp 0
transform 1 0 17986 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_43_333
timestamp 0
transform 1 0 18354 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_43_346
timestamp 0
transform 1 0 18952 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_43_354
timestamp 0
transform 1 0 19320 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_43_358
timestamp 0
transform 1 0 19504 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_43_361
timestamp 0
transform 1 0 19642 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_369
timestamp 0
transform 1 0 20010 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_43_377
timestamp 0
transform 1 0 20378 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_379
timestamp 0
transform 1 0 20470 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_43_404
timestamp 0
transform 1 0 21620 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_412
timestamp 0
transform 1 0 21988 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_421
timestamp 0
transform 1 0 22402 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_429
timestamp 0
transform 1 0 22770 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_437
timestamp 0
transform 1 0 23138 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_445
timestamp 0
transform 1 0 23506 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_453
timestamp 0
transform 1 0 23874 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_461
timestamp 0
transform 1 0 24242 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_469
timestamp 0
transform 1 0 24610 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_43_477
timestamp 0
transform 1 0 24978 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_479
timestamp 0
transform 1 0 25070 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_43_481
timestamp 0
transform 1 0 25162 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_489
timestamp 0
transform 1 0 25530 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_497
timestamp 0
transform 1 0 25898 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_505
timestamp 0
transform 1 0 26266 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_513
timestamp 0
transform 1 0 26634 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_521
timestamp 0
transform 1 0 27002 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_43_529
timestamp 0
transform 1 0 27370 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_43_537
timestamp 0
transform 1 0 27738 0 -1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_43_539
timestamp 0
transform 1 0 27830 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_43_541
timestamp 0
transform 1 0 27922 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_43_549
timestamp 0
transform 1 0 28290 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_43_574
timestamp 0
transform 1 0 29440 0 -1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_43_582
timestamp 0
transform 1 0 29808 0 -1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_44_0
timestamp 0
transform 1 0 3036 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_8
timestamp 0
transform 1 0 3404 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_16
timestamp 0
transform 1 0 3772 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_24
timestamp 0
transform 1 0 4140 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_44_28
timestamp 0
transform 1 0 4324 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_44_31
timestamp 0
transform 1 0 4462 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_39
timestamp 0
transform 1 0 4830 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_47
timestamp 0
transform 1 0 5198 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_79
timestamp 0
transform 1 0 6670 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_44_87
timestamp 0
transform 1 0 7038 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 0
transform 1 0 7130 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_91
timestamp 0
transform 1 0 7222 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_99
timestamp 0
transform 1 0 7590 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_44_103
timestamp 0
transform 1 0 7774 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_128
timestamp 0
transform 1 0 8924 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_136
timestamp 0
transform 1 0 9292 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_144
timestamp 0
transform 1 0 9660 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_44_148
timestamp 0
transform 1 0 9844 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_44_151
timestamp 0
transform 1 0 9982 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_159
timestamp 0
transform 1 0 10350 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_44_167
timestamp 0
transform 1 0 10718 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_44_169
timestamp 0
transform 1 0 10810 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_194
timestamp 0
transform 1 0 11960 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_202
timestamp 0
transform 1 0 12328 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_211
timestamp 0
transform 1 0 12742 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_219
timestamp 0
transform 1 0 13110 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_227
timestamp 0
transform 1 0 13478 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_44_231
timestamp 0
transform 1 0 13662 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_44_233
timestamp 0
transform 1 0 13754 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_258
timestamp 0
transform 1 0 14904 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_266
timestamp 0
transform 1 0 15272 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_44_271
timestamp 0
transform 1 0 15502 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_44_275
timestamp 0
transform 1 0 15686 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_44_283
timestamp 0
transform 1 0 16054 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_44_293
timestamp 0
transform 1 0 16514 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_44_301
timestamp 0
transform 1 0 16882 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_44_326
timestamp 0
transform 1 0 18032 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_44_331
timestamp 0
transform 1 0 18262 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_44_359
timestamp 0
transform 1 0 19550 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_44_367
timestamp 0
transform 1 0 19918 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_374
timestamp 0
transform 1 0 20240 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_382
timestamp 0
transform 1 0 20608 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_391
timestamp 0
transform 1 0 21022 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_399
timestamp 0
transform 1 0 21390 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_407
timestamp 0
transform 1 0 21758 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_415
timestamp 0
transform 1 0 22126 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_423
timestamp 0
transform 1 0 22494 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_44_427
timestamp 0
transform 1 0 22678 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_433
timestamp 0
transform 1 0 22954 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_441
timestamp 0
transform 1 0 23322 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_44_449
timestamp 0
transform 1 0 23690 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_451
timestamp 0
transform 1 0 23782 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_44_459
timestamp 0
transform 1 0 24150 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_44_485
timestamp 0
transform 1 0 25346 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_493
timestamp 0
transform 1 0 25714 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_501
timestamp 0
transform 1 0 26082 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_44_509
timestamp 0
transform 1 0 26450 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_44_511
timestamp 0
transform 1 0 26542 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_44_539
timestamp 0
transform 1 0 27830 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_547
timestamp 0
transform 1 0 28198 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_44_555
timestamp 0
transform 1 0 28566 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_563
timestamp 0
transform 1 0 28934 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_44_567
timestamp 0
transform 1 0 29118 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_44_569
timestamp 0
transform 1 0 29210 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_44_571
timestamp 0
transform 1 0 29302 0 1 15232
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_44_579
timestamp 0
transform 1 0 29670 0 1 15232
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_44_583
timestamp 0
transform 1 0 29854 0 1 15232
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_44_585
timestamp 0
transform 1 0 29946 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_0
timestamp 0
transform 1 0 3036 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_45_8
timestamp 0
transform 1 0 3404 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_33
timestamp 0
transform 1 0 4554 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_41
timestamp 0
transform 1 0 4922 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_49
timestamp 0
transform 1 0 5290 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 0
transform 1 0 5658 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_45_59
timestamp 0
transform 1 0 5750 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_61
timestamp 0
transform 1 0 5842 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_69
timestamp 0
transform 1 0 6210 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_77
timestamp 0
transform 1 0 6578 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_85
timestamp 0
transform 1 0 6946 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_93
timestamp 0
transform 1 0 7314 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_101
timestamp 0
transform 1 0 7682 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_109
timestamp 0
transform 1 0 8050 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_45_117
timestamp 0
transform 1 0 8418 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_45_119
timestamp 0
transform 1 0 8510 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_121
timestamp 0
transform 1 0 8602 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_45_129
timestamp 0
transform 1 0 8970 0 -1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_45_133
timestamp 0
transform 1 0 9154 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_158
timestamp 0
transform 1 0 10304 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_166
timestamp 0
transform 1 0 10672 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_45_174
timestamp 0
transform 1 0 11040 0 -1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_45_178
timestamp 0
transform 1 0 11224 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_45_181
timestamp 0
transform 1 0 11362 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_189
timestamp 0
transform 1 0 11730 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_197
timestamp 0
transform 1 0 12098 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_229
timestamp 0
transform 1 0 13570 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_45_237
timestamp 0
transform 1 0 13938 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 0
transform 1 0 14030 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_241
timestamp 0
transform 1 0 14122 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_249
timestamp 0
transform 1 0 14490 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_257
timestamp 0
transform 1 0 14858 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_45_265
timestamp 0
transform 1 0 15226 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_45_291
timestamp 0
transform 1 0 16422 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_45_299
timestamp 0
transform 1 0 16790 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_301
timestamp 0
transform 1 0 16882 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_309
timestamp 0
transform 1 0 17250 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_317
timestamp 0
transform 1 0 17618 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_45_325
timestamp 0
transform 1 0 17986 0 -1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_45_329
timestamp 0
transform 1 0 18170 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_45_331
timestamp 0
transform 1 0 18262 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_45_356
timestamp 0
transform 1 0 19412 0 -1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_45_361
timestamp 0
transform 1 0 19642 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_45_369
timestamp 0
transform 1 0 20010 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_394
timestamp 0
transform 1 0 21160 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_45_402
timestamp 0
transform 1 0 21528 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_411
timestamp 0
transform 1 0 21942 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_45_419
timestamp 0
transform 1 0 22310 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_421
timestamp 0
transform 1 0 22402 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_429
timestamp 0
transform 1 0 22770 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_437
timestamp 0
transform 1 0 23138 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_445
timestamp 0
transform 1 0 23506 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_453
timestamp 0
transform 1 0 23874 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_461
timestamp 0
transform 1 0 24242 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_469
timestamp 0
transform 1 0 24610 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_45_477
timestamp 0
transform 1 0 24978 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_45_479
timestamp 0
transform 1 0 25070 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_45_481
timestamp 0
transform 1 0 25162 0 -1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_45_509
timestamp 0
transform 1 0 26450 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_45_517
timestamp 0
transform 1 0 26818 0 -1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_45_521
timestamp 0
transform 1 0 27002 0 -1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_45_523
timestamp 0
transform 1 0 27094 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_45_532
timestamp 0
transform 1 0 27508 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_541
timestamp 0
transform 1 0 27922 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_549
timestamp 0
transform 1 0 28290 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_557
timestamp 0
transform 1 0 28658 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_565
timestamp 0
transform 1 0 29026 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_45_573
timestamp 0
transform 1 0 29394 0 -1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_45_581
timestamp 0
transform 1 0 29762 0 -1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_45_585
timestamp 0
transform 1 0 29946 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_46_0
timestamp 0
transform 1 0 3036 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_46_26
timestamp 0
transform 1 0 4232 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_46_31
timestamp 0
transform 1 0 4462 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_46_39
timestamp 0
transform 1 0 4830 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_46_43
timestamp 0
transform 1 0 5014 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_45
timestamp 0
transform 1 0 5106 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_46_70
timestamp 0
transform 1 0 6256 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_78
timestamp 0
transform 1 0 6624 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_46_86
timestamp 0
transform 1 0 6992 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_46_91
timestamp 0
transform 1 0 7222 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_99
timestamp 0
transform 1 0 7590 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_107
timestamp 0
transform 1 0 7958 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_109
timestamp 0
transform 1 0 8050 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_46_118
timestamp 0
transform 1 0 8464 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_126
timestamp 0
transform 1 0 8832 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_134
timestamp 0
transform 1 0 9200 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_142
timestamp 0
transform 1 0 9568 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_151
timestamp 0
transform 1 0 9982 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_159
timestamp 0
transform 1 0 10350 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_46_167
timestamp 0
transform 1 0 10718 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_46_192
timestamp 0
transform 1 0 11868 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_200
timestamp 0
transform 1 0 12236 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_208
timestamp 0
transform 1 0 12604 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_46_211
timestamp 0
transform 1 0 12742 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_219
timestamp 0
transform 1 0 13110 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_227
timestamp 0
transform 1 0 13478 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_235
timestamp 0
transform 1 0 13846 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_243
timestamp 0
transform 1 0 14214 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_251
timestamp 0
transform 1 0 14582 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_259
timestamp 0
transform 1 0 14950 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_267
timestamp 0
transform 1 0 15318 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_269
timestamp 0
transform 1 0 15410 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_46_271
timestamp 0
transform 1 0 15502 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_279
timestamp 0
transform 1 0 15870 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_287
timestamp 0
transform 1 0 16238 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_295
timestamp 0
transform 1 0 16606 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_303
timestamp 0
transform 1 0 16974 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_311
timestamp 0
transform 1 0 17342 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_319
timestamp 0
transform 1 0 17710 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_327
timestamp 0
transform 1 0 18078 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_329
timestamp 0
transform 1 0 18170 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_46_331
timestamp 0
transform 1 0 18262 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_339
timestamp 0
transform 1 0 18630 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_347
timestamp 0
transform 1 0 18998 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_355
timestamp 0
transform 1 0 19366 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_363
timestamp 0
transform 1 0 19734 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_371
timestamp 0
transform 1 0 20102 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_379
timestamp 0
transform 1 0 20470 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_387
timestamp 0
transform 1 0 20838 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_389
timestamp 0
transform 1 0 20930 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_46_391
timestamp 0
transform 1 0 21022 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_399
timestamp 0
transform 1 0 21390 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_407
timestamp 0
transform 1 0 21758 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_415
timestamp 0
transform 1 0 22126 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_423
timestamp 0
transform 1 0 22494 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_431
timestamp 0
transform 1 0 22862 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_439
timestamp 0
transform 1 0 23230 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_447
timestamp 0
transform 1 0 23598 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_449
timestamp 0
transform 1 0 23690 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_46_451
timestamp 0
transform 1 0 23782 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_46_459
timestamp 0
transform 1 0 24150 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_46_487
timestamp 0
transform 1 0 25438 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_46_499
timestamp 0
transform 1 0 25990 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_507
timestamp 0
transform 1 0 26358 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_509
timestamp 0
transform 1 0 26450 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_46_511
timestamp 0
transform 1 0 26542 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_46_539
timestamp 0
transform 1 0 27830 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_46_547
timestamp 0
transform 1 0 28198 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_46_555
timestamp 0
transform 1 0 28566 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_557
timestamp 0
transform 1 0 28658 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_46_566
timestamp 0
transform 1 0 29072 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_46_571
timestamp 0
transform 1 0 29302 0 1 15776
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_46_579
timestamp 0
transform 1 0 29670 0 1 15776
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_46_583
timestamp 0
transform 1 0 29854 0 1 15776
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_46_585
timestamp 0
transform 1 0 29946 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_47_0
timestamp 0
transform 1 0 3036 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_47_28
timestamp 0
transform 1 0 4324 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_47_56
timestamp 0
transform 1 0 5612 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_47_61
timestamp 0
transform 1 0 5842 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_47_65
timestamp 0
transform 1 0 6026 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_47_74
timestamp 0
transform 1 0 6440 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_47_82
timestamp 0
transform 1 0 6808 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_47_90
timestamp 0
transform 1 0 7176 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_47_115
timestamp 0
transform 1 0 8326 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_47_119
timestamp 0
transform 1 0 8510 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_47_121
timestamp 0
transform 1 0 8602 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_47_149
timestamp 0
transform 1 0 9890 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_157
timestamp 0
transform 1 0 10258 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_165
timestamp 0
transform 1 0 10626 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_47_173
timestamp 0
transform 1 0 10994 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_47_177
timestamp 0
transform 1 0 11178 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_47_179
timestamp 0
transform 1 0 11270 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_47_181
timestamp 0
transform 1 0 11362 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_189
timestamp 0
transform 1 0 11730 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_197
timestamp 0
transform 1 0 12098 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_47_205
timestamp 0
transform 1 0 12466 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_47_209
timestamp 0
transform 1 0 12650 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_47_234
timestamp 0
transform 1 0 13800 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_47_238
timestamp 0
transform 1 0 13984 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_47_241
timestamp 0
transform 1 0 14122 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_249
timestamp 0
transform 1 0 14490 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_257
timestamp 0
transform 1 0 14858 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_265
timestamp 0
transform 1 0 15226 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_273
timestamp 0
transform 1 0 15594 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_281
timestamp 0
transform 1 0 15962 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_289
timestamp 0
transform 1 0 16330 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_47_297
timestamp 0
transform 1 0 16698 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_47_299
timestamp 0
transform 1 0 16790 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_47_301
timestamp 0
transform 1 0 16882 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_309
timestamp 0
transform 1 0 17250 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_317
timestamp 0
transform 1 0 17618 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_325
timestamp 0
transform 1 0 17986 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_333
timestamp 0
transform 1 0 18354 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_341
timestamp 0
transform 1 0 18722 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_349
timestamp 0
transform 1 0 19090 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_47_357
timestamp 0
transform 1 0 19458 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_47_359
timestamp 0
transform 1 0 19550 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_47_361
timestamp 0
transform 1 0 19642 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_369
timestamp 0
transform 1 0 20010 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_377
timestamp 0
transform 1 0 20378 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_409
timestamp 0
transform 1 0 21850 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_47_417
timestamp 0
transform 1 0 22218 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_47_419
timestamp 0
transform 1 0 22310 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_47_421
timestamp 0
transform 1 0 22402 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_47_429
timestamp 0
transform 1 0 22770 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_47_454
timestamp 0
transform 1 0 23920 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_462
timestamp 0
transform 1 0 24288 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_470
timestamp 0
transform 1 0 24656 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_47_478
timestamp 0
transform 1 0 25024 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_47_481
timestamp 0
transform 1 0 25162 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_489
timestamp 0
transform 1 0 25530 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_521
timestamp 0
transform 1 0 27002 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_529
timestamp 0
transform 1 0 27370 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_47_537
timestamp 0
transform 1 0 27738 0 -1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_47_539
timestamp 0
transform 1 0 27830 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_47_541
timestamp 0
transform 1 0 27922 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_47_573
timestamp 0
transform 1 0 29394 0 -1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_47_581
timestamp 0
transform 1 0 29762 0 -1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_47_585
timestamp 0
transform 1 0 29946 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_48_0
timestamp 0
transform 1 0 3036 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_8
timestamp 0
transform 1 0 3404 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_16
timestamp 0
transform 1 0 3772 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_48_24
timestamp 0
transform 1 0 4140 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_48_28
timestamp 0
transform 1 0 4324 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_48_31
timestamp 0
transform 1 0 4462 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_48_43
timestamp 0
transform 1 0 5014 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_48_51
timestamp 0
transform 1 0 5382 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_48_55
timestamp 0
transform 1 0 5566 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_48_57
timestamp 0
transform 1 0 5658 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_48_82
timestamp 0
transform 1 0 6808 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_48_91
timestamp 0
transform 1 0 7222 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_48_111
timestamp 0
transform 1 0 8142 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_48_119
timestamp 0
transform 1 0 8510 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_48_121
timestamp 0
transform 1 0 8602 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_48_146
timestamp 0
transform 1 0 9752 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_48_151
timestamp 0
transform 1 0 9982 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_48_159
timestamp 0
transform 1 0 10350 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_48_163
timestamp 0
transform 1 0 10534 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_48_188
timestamp 0
transform 1 0 11684 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_196
timestamp 0
transform 1 0 12052 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_48_204
timestamp 0
transform 1 0 12420 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_48_208
timestamp 0
transform 1 0 12604 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_48_211
timestamp 0
transform 1 0 12742 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_219
timestamp 0
transform 1 0 13110 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_48_227
timestamp 0
transform 1 0 13478 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_48_231
timestamp 0
transform 1 0 13662 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_48_233
timestamp 0
transform 1 0 13754 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_48_258
timestamp 0
transform 1 0 14904 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_48_266
timestamp 0
transform 1 0 15272 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_48_271
timestamp 0
transform 1 0 15502 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_48_279
timestamp 0
transform 1 0 15870 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_48_304
timestamp 0
transform 1 0 17020 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_48_311
timestamp 0
transform 1 0 17342 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_319
timestamp 0
transform 1 0 17710 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_48_327
timestamp 0
transform 1 0 18078 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_48_329
timestamp 0
transform 1 0 18170 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_48_331
timestamp 0
transform 1 0 18262 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_339
timestamp 0
transform 1 0 18630 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_347
timestamp 0
transform 1 0 18998 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_355
timestamp 0
transform 1 0 19366 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_363
timestamp 0
transform 1 0 19734 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_371
timestamp 0
transform 1 0 20102 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_379
timestamp 0
transform 1 0 20470 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_48_387
timestamp 0
transform 1 0 20838 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_48_389
timestamp 0
transform 1 0 20930 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_48_391
timestamp 0
transform 1 0 21022 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_399
timestamp 0
transform 1 0 21390 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_407
timestamp 0
transform 1 0 21758 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_415
timestamp 0
transform 1 0 22126 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_423
timestamp 0
transform 1 0 22494 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_431
timestamp 0
transform 1 0 22862 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_439
timestamp 0
transform 1 0 23230 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_48_447
timestamp 0
transform 1 0 23598 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_48_449
timestamp 0
transform 1 0 23690 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_48_451
timestamp 0
transform 1 0 23782 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_48_461
timestamp 0
transform 1 0 24242 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_469
timestamp 0
transform 1 0 24610 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_477
timestamp 0
transform 1 0 24978 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_485
timestamp 0
transform 1 0 25346 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_493
timestamp 0
transform 1 0 25714 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_501
timestamp 0
transform 1 0 26082 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_48_509
timestamp 0
transform 1 0 26450 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_48_511
timestamp 0
transform 1 0 26542 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_519
timestamp 0
transform 1 0 26910 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_527
timestamp 0
transform 1 0 27278 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_535
timestamp 0
transform 1 0 27646 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_543
timestamp 0
transform 1 0 28014 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_551
timestamp 0
transform 1 0 28382 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_48_559
timestamp 0
transform 1 0 28750 0 1 16320
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_48_567
timestamp 0
transform 1 0 29118 0 1 16320
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_48_569
timestamp 0
transform 1 0 29210 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_48_571
timestamp 0
transform 1 0 29302 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_48_581
timestamp 0
transform 1 0 29762 0 1 16320
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_48_585
timestamp 0
transform 1 0 29946 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_49_0
timestamp 0
transform 1 0 3036 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_8
timestamp 0
transform 1 0 3404 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_16
timestamp 0
transform 1 0 3772 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_24
timestamp 0
transform 1 0 4140 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_32
timestamp 0
transform 1 0 4508 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_40
timestamp 0
transform 1 0 4876 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_48
timestamp 0
transform 1 0 5244 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_56
timestamp 0
transform 1 0 5612 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_49_61
timestamp 0
transform 1 0 5842 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_69
timestamp 0
transform 1 0 6210 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_77
timestamp 0
transform 1 0 6578 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_85
timestamp 0
transform 1 0 6946 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 0
transform 1 0 7130 0 -1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_49_91
timestamp 0
transform 1 0 7222 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_49_116
timestamp 0
transform 1 0 8372 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_49_121
timestamp 0
transform 1 0 8602 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_129
timestamp 0
transform 1 0 8970 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_137
timestamp 0
transform 1 0 9338 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_49_148
timestamp 0
transform 1 0 9844 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_49_176
timestamp 0
transform 1 0 11132 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_49_181
timestamp 0
transform 1 0 11362 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_49_191
timestamp 0
transform 1 0 11822 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_49_198
timestamp 0
transform 1 0 12144 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_206
timestamp 0
transform 1 0 12512 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_49_210
timestamp 0
transform 1 0 12696 0 -1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_49_236
timestamp 0
transform 1 0 13892 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_49_241
timestamp 0
transform 1 0 14122 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_49_253
timestamp 0
transform 1 0 14674 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_49_264
timestamp 0
transform 1 0 15180 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_296
timestamp 0
transform 1 0 16652 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_49_301
timestamp 0
transform 1 0 16882 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_49_311
timestamp 0
transform 1 0 17342 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_49_319
timestamp 0
transform 1 0 17710 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_49_344
timestamp 0
transform 1 0 18860 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_352
timestamp 0
transform 1 0 19228 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_361
timestamp 0
transform 1 0 19642 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_393
timestamp 0
transform 1 0 21114 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_49_405
timestamp 0
transform 1 0 21666 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_413
timestamp 0
transform 1 0 22034 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_49_417
timestamp 0
transform 1 0 22218 0 -1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_49_419
timestamp 0
transform 1 0 22310 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_49_421
timestamp 0
transform 1 0 22402 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_429
timestamp 0
transform 1 0 22770 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_49_457
timestamp 0
transform 1 0 24058 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_465
timestamp 0
transform 1 0 24426 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_49_473
timestamp 0
transform 1 0 24794 0 -1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_49_477
timestamp 0
transform 1 0 24978 0 -1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_49_479
timestamp 0
transform 1 0 25070 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_49_481
timestamp 0
transform 1 0 25162 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_489
timestamp 0
transform 1 0 25530 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_49_497
timestamp 0
transform 1 0 25898 0 -1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_49_523
timestamp 0
transform 1 0 27094 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_49_531
timestamp 0
transform 1 0 27462 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_49_539
timestamp 0
transform 1 0 27830 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_49_541
timestamp 0
transform 1 0 27922 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_49_549
timestamp 0
transform 1 0 28290 0 -1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_49_575
timestamp 0
transform 1 0 29486 0 -1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_49_583
timestamp 0
transform 1 0 29854 0 -1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_49_585
timestamp 0
transform 1 0 29946 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_50_0
timestamp 0
transform 1 0 3036 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_8
timestamp 0
transform 1 0 3404 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_16
timestamp 0
transform 1 0 3772 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_24
timestamp 0
transform 1 0 4140 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_28
timestamp 0
transform 1 0 4324 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_50_31
timestamp 0
transform 1 0 4462 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_39
timestamp 0
transform 1 0 4830 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_47
timestamp 0
transform 1 0 5198 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_51
timestamp 0
transform 1 0 5382 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_50_77
timestamp 0
transform 1 0 6578 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_85
timestamp 0
transform 1 0 6946 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 0
transform 1 0 7130 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_50_91
timestamp 0
transform 1 0 7222 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_99
timestamp 0
transform 1 0 7590 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_107
timestamp 0
transform 1 0 7958 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_115
timestamp 0
transform 1 0 8326 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_119
timestamp 0
transform 1 0 8510 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 0
transform 1 0 8602 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_146
timestamp 0
transform 1 0 9752 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_50_151
timestamp 0
transform 1 0 9982 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_159
timestamp 0
transform 1 0 10350 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_167
timestamp 0
transform 1 0 10718 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_50_171
timestamp 0
transform 1 0 10902 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_196
timestamp 0
transform 1 0 12052 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_50_203
timestamp 0
transform 1 0 12374 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_207
timestamp 0
transform 1 0 12558 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_50_209
timestamp 0
transform 1 0 12650 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_211
timestamp 0
transform 1 0 12742 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_50_239
timestamp 0
transform 1 0 14030 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_247
timestamp 0
transform 1 0 14398 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 0
transform 1 0 14582 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_258
timestamp 0
transform 1 0 14904 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_50_262
timestamp 0
transform 1 0 15088 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_266
timestamp 0
transform 1 0 15272 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_50_271
timestamp 0
transform 1 0 15502 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_275
timestamp 0
transform 1 0 15686 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_50_301
timestamp 0
transform 1 0 16882 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_50_308
timestamp 0
transform 1 0 17204 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_316
timestamp 0
transform 1 0 17572 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_324
timestamp 0
transform 1 0 17940 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_328
timestamp 0
transform 1 0 18124 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_50_331
timestamp 0
transform 1 0 18262 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_339
timestamp 0
transform 1 0 18630 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_347
timestamp 0
transform 1 0 18998 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_355
timestamp 0
transform 1 0 19366 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_363
timestamp 0
transform 1 0 19734 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_371
timestamp 0
transform 1 0 20102 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_379
timestamp 0
transform 1 0 20470 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_50_387
timestamp 0
transform 1 0 20838 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_50_389
timestamp 0
transform 1 0 20930 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_391
timestamp 0
transform 1 0 21022 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_50_419
timestamp 0
transform 1 0 22310 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_427
timestamp 0
transform 1 0 22678 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_435
timestamp 0
transform 1 0 23046 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_443
timestamp 0
transform 1 0 23414 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_447
timestamp 0
transform 1 0 23598 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_50_449
timestamp 0
transform 1 0 23690 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_50_451
timestamp 0
transform 1 0 23782 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_459
timestamp 0
transform 1 0 24150 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_491
timestamp 0
transform 1 0 25622 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_499
timestamp 0
transform 1 0 25990 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_50_507
timestamp 0
transform 1 0 26358 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_50_509
timestamp 0
transform 1 0 26450 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_511
timestamp 0
transform 1 0 26542 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_50_539
timestamp 0
transform 1 0 27830 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_50_547
timestamp 0
transform 1 0 28198 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_50_555
timestamp 0
transform 1 0 28566 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_50_565
timestamp 0
transform 1 0 29026 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_50_569
timestamp 0
transform 1 0 29210 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_50_571
timestamp 0
transform 1 0 29302 0 1 16864
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_50_579
timestamp 0
transform 1 0 29670 0 1 16864
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_50_583
timestamp 0
transform 1 0 29854 0 1 16864
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_50_585
timestamp 0
transform 1 0 29946 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_51_0
timestamp 0
transform 1 0 3036 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_8
timestamp 0
transform 1 0 3404 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_51_36
timestamp 0
transform 1 0 4692 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_44
timestamp 0
transform 1 0 5060 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_52
timestamp 0
transform 1 0 5428 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_61
timestamp 0
transform 1 0 5842 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_69
timestamp 0
transform 1 0 6210 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_77
timestamp 0
transform 1 0 6578 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_85
timestamp 0
transform 1 0 6946 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_51_89
timestamp 0
transform 1 0 7130 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_51_115
timestamp 0
transform 1 0 8326 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_51_119
timestamp 0
transform 1 0 8510 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_51_121
timestamp 0
transform 1 0 8602 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_129
timestamp 0
transform 1 0 8970 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_137
timestamp 0
transform 1 0 9338 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_145
timestamp 0
transform 1 0 9706 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_153
timestamp 0
transform 1 0 10074 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_161
timestamp 0
transform 1 0 10442 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_169
timestamp 0
transform 1 0 10810 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_51_177
timestamp 0
transform 1 0 11178 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_51_179
timestamp 0
transform 1 0 11270 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_51_181
timestamp 0
transform 1 0 11362 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_189
timestamp 0
transform 1 0 11730 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_197
timestamp 0
transform 1 0 12098 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_51_205
timestamp 0
transform 1 0 12466 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_51_207
timestamp 0
transform 1 0 12558 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_51_232
timestamp 0
transform 1 0 13708 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_241
timestamp 0
transform 1 0 14122 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_249
timestamp 0
transform 1 0 14490 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_51_277
timestamp 0
transform 1 0 15778 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_285
timestamp 0
transform 1 0 16146 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_293
timestamp 0
transform 1 0 16514 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 0
transform 1 0 16698 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_51_299
timestamp 0
transform 1 0 16790 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_51_301
timestamp 0
transform 1 0 16882 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_309
timestamp 0
transform 1 0 17250 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_51_317
timestamp 0
transform 1 0 17618 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_51_343
timestamp 0
transform 1 0 18814 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_351
timestamp 0
transform 1 0 19182 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_51_359
timestamp 0
transform 1 0 19550 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_51_361
timestamp 0
transform 1 0 19642 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_369
timestamp 0
transform 1 0 20010 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_51_373
timestamp 0
transform 1 0 20194 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_51_398
timestamp 0
transform 1 0 21344 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_406
timestamp 0
transform 1 0 21712 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_414
timestamp 0
transform 1 0 22080 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_51_418
timestamp 0
transform 1 0 22264 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_51_421
timestamp 0
transform 1 0 22402 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_429
timestamp 0
transform 1 0 22770 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_51_457
timestamp 0
transform 1 0 24058 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_51_465
timestamp 0
transform 1 0 24426 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_473
timestamp 0
transform 1 0 24794 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_51_477
timestamp 0
transform 1 0 24978 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_51_479
timestamp 0
transform 1 0 25070 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_51_481
timestamp 0
transform 1 0 25162 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_51_509
timestamp 0
transform 1 0 26450 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_51_517
timestamp 0
transform 1 0 26818 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_51_521
timestamp 0
transform 1 0 27002 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_51_531
timestamp 0
transform 1 0 27462 0 -1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_51_539
timestamp 0
transform 1 0 27830 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_51_541
timestamp 0
transform 1 0 27922 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_51_545
timestamp 0
transform 1 0 28106 0 -1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_51_571
timestamp 0
transform 1 0 29302 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_51_581
timestamp 0
transform 1 0 29762 0 -1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_51_585
timestamp 0
transform 1 0 29946 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_52_0
timestamp 0
transform 1 0 3036 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_52_26
timestamp 0
transform 1 0 4232 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_52_31
timestamp 0
transform 1 0 4462 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_52_41
timestamp 0
transform 1 0 4922 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_52_49
timestamp 0
transform 1 0 5290 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_52_53
timestamp 0
transform 1 0 5474 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_55
timestamp 0
transform 1 0 5566 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_52_80
timestamp 0
transform 1 0 6716 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_52_88
timestamp 0
transform 1 0 7084 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_52_91
timestamp 0
transform 1 0 7222 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_99
timestamp 0
transform 1 0 7590 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_52_107
timestamp 0
transform 1 0 7958 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_52_111
timestamp 0
transform 1 0 8142 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_52_137
timestamp 0
transform 1 0 9338 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_52_145
timestamp 0
transform 1 0 9706 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_52_149
timestamp 0
transform 1 0 9890 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_52_151
timestamp 0
transform 1 0 9982 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_159
timestamp 0
transform 1 0 10350 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_167
timestamp 0
transform 1 0 10718 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_175
timestamp 0
transform 1 0 11086 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_183
timestamp 0
transform 1 0 11454 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_191
timestamp 0
transform 1 0 11822 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_199
timestamp 0
transform 1 0 12190 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_52_207
timestamp 0
transform 1 0 12558 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_209
timestamp 0
transform 1 0 12650 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_52_211
timestamp 0
transform 1 0 12742 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_219
timestamp 0
transform 1 0 13110 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_227
timestamp 0
transform 1 0 13478 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_235
timestamp 0
transform 1 0 13846 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_243
timestamp 0
transform 1 0 14214 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_251
timestamp 0
transform 1 0 14582 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_259
timestamp 0
transform 1 0 14950 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_52_267
timestamp 0
transform 1 0 15318 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_269
timestamp 0
transform 1 0 15410 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_52_271
timestamp 0
transform 1 0 15502 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_279
timestamp 0
transform 1 0 15870 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_287
timestamp 0
transform 1 0 16238 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_295
timestamp 0
transform 1 0 16606 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_303
timestamp 0
transform 1 0 16974 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_311
timestamp 0
transform 1 0 17342 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_319
timestamp 0
transform 1 0 17710 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_52_327
timestamp 0
transform 1 0 18078 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_329
timestamp 0
transform 1 0 18170 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_52_331
timestamp 0
transform 1 0 18262 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_52_339
timestamp 0
transform 1 0 18630 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_341
timestamp 0
transform 1 0 18722 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_52_350
timestamp 0
transform 1 0 19136 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_358
timestamp 0
transform 1 0 19504 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_366
timestamp 0
transform 1 0 19872 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_374
timestamp 0
transform 1 0 20240 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_382
timestamp 0
transform 1 0 20608 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_391
timestamp 0
transform 1 0 21022 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_399
timestamp 0
transform 1 0 21390 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_407
timestamp 0
transform 1 0 21758 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_52_415
timestamp 0
transform 1 0 22126 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_52_419
timestamp 0
transform 1 0 22310 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_421
timestamp 0
transform 1 0 22402 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_52_446
timestamp 0
transform 1 0 23552 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_52_451
timestamp 0
transform 1 0 23782 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_52_459
timestamp 0
transform 1 0 24150 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_52_463
timestamp 0
transform 1 0 24334 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_465
timestamp 0
transform 1 0 24426 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_52_490
timestamp 0
transform 1 0 25576 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_52_502
timestamp 0
transform 1 0 26128 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_511
timestamp 0
transform 1 0 26542 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_519
timestamp 0
transform 1 0 26910 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_52_527
timestamp 0
transform 1 0 27278 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_52_535
timestamp 0
transform 1 0 27646 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_52_539
timestamp 0
transform 1 0 27830 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_541
timestamp 0
transform 1 0 27922 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_52_566
timestamp 0
transform 1 0 29072 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_52_571
timestamp 0
transform 1 0 29302 0 1 17408
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_52_579
timestamp 0
transform 1 0 29670 0 1 17408
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_52_583
timestamp 0
transform 1 0 29854 0 1 17408
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_52_585
timestamp 0
transform 1 0 29946 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_53_0
timestamp 0
transform 1 0 3036 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_8
timestamp 0
transform 1 0 3404 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_16
timestamp 0
transform 1 0 3772 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_24
timestamp 0
transform 1 0 4140 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_32
timestamp 0
transform 1 0 4508 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_40
timestamp 0
transform 1 0 4876 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_48
timestamp 0
transform 1 0 5244 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_53_56
timestamp 0
transform 1 0 5612 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_53_61
timestamp 0
transform 1 0 5842 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_69
timestamp 0
transform 1 0 6210 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_53_77
timestamp 0
transform 1 0 6578 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_53_103
timestamp 0
transform 1 0 7774 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_111
timestamp 0
transform 1 0 8142 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_53_119
timestamp 0
transform 1 0 8510 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_53_121
timestamp 0
transform 1 0 8602 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_129
timestamp 0
transform 1 0 8970 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_137
timestamp 0
transform 1 0 9338 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_145
timestamp 0
transform 1 0 9706 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_153
timestamp 0
transform 1 0 10074 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_161
timestamp 0
transform 1 0 10442 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_169
timestamp 0
transform 1 0 10810 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_53_177
timestamp 0
transform 1 0 11178 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_53_179
timestamp 0
transform 1 0 11270 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_53_181
timestamp 0
transform 1 0 11362 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_189
timestamp 0
transform 1 0 11730 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_197
timestamp 0
transform 1 0 12098 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_53_205
timestamp 0
transform 1 0 12466 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_53_209
timestamp 0
transform 1 0 12650 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_53_211
timestamp 0
transform 1 0 12742 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_53_236
timestamp 0
transform 1 0 13892 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_53_241
timestamp 0
transform 1 0 14122 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_249
timestamp 0
transform 1 0 14490 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_257
timestamp 0
transform 1 0 14858 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_265
timestamp 0
transform 1 0 15226 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_273
timestamp 0
transform 1 0 15594 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_281
timestamp 0
transform 1 0 15962 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_289
timestamp 0
transform 1 0 16330 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 0
transform 1 0 16698 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_53_299
timestamp 0
transform 1 0 16790 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_53_301
timestamp 0
transform 1 0 16882 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_309
timestamp 0
transform 1 0 17250 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_317
timestamp 0
transform 1 0 17618 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_325
timestamp 0
transform 1 0 17986 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_333
timestamp 0
transform 1 0 18354 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_53_341
timestamp 0
transform 1 0 18722 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_53_345
timestamp 0
transform 1 0 18906 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_53_353
timestamp 0
transform 1 0 19274 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_53_357
timestamp 0
transform 1 0 19458 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_53_359
timestamp 0
transform 1 0 19550 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_53_361
timestamp 0
transform 1 0 19642 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_369
timestamp 0
transform 1 0 20010 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_377
timestamp 0
transform 1 0 20378 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_53_385
timestamp 0
transform 1 0 20746 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_53_389
timestamp 0
transform 1 0 20930 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 0
transform 1 0 21022 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_53_416
timestamp 0
transform 1 0 22172 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_53_421
timestamp 0
transform 1 0 22402 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_53_425
timestamp 0
transform 1 0 22586 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_53_427
timestamp 0
transform 1 0 22678 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_53_452
timestamp 0
transform 1 0 23828 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_53_464
timestamp 0
transform 1 0 24380 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_472
timestamp 0
transform 1 0 24748 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_481
timestamp 0
transform 1 0 25162 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_489
timestamp 0
transform 1 0 25530 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_53_497
timestamp 0
transform 1 0 25898 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_53_501
timestamp 0
transform 1 0 26082 0 -1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 0
transform 1 0 26174 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_53_528
timestamp 0
transform 1 0 27324 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_53_536
timestamp 0
transform 1 0 27692 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_53_541
timestamp 0
transform 1 0 27922 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_549
timestamp 0
transform 1 0 28290 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_557
timestamp 0
transform 1 0 28658 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_565
timestamp 0
transform 1 0 29026 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_53_573
timestamp 0
transform 1 0 29394 0 -1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_53_581
timestamp 0
transform 1 0 29762 0 -1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_53_585
timestamp 0
transform 1 0 29946 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_54_0
timestamp 0
transform 1 0 3036 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_54_26
timestamp 0
transform 1 0 4232 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_54_31
timestamp 0
transform 1 0 4462 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_39
timestamp 0
transform 1 0 4830 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_54_43
timestamp 0
transform 1 0 5014 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_45
timestamp 0
transform 1 0 5106 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_66
timestamp 0
transform 1 0 6072 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_74
timestamp 0
transform 1 0 6440 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_54_78
timestamp 0
transform 1 0 6624 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_54_86
timestamp 0
transform 1 0 6992 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_54_91
timestamp 0
transform 1 0 7222 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_54_102
timestamp 0
transform 1 0 7728 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_110
timestamp 0
transform 1 0 8096 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_54_114
timestamp 0
transform 1 0 8280 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_116
timestamp 0
transform 1 0 8372 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_141
timestamp 0
transform 1 0 9522 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_54_149
timestamp 0
transform 1 0 9890 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_54_151
timestamp 0
transform 1 0 9982 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_54_179
timestamp 0
transform 1 0 11270 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_187
timestamp 0
transform 1 0 11638 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_195
timestamp 0
transform 1 0 12006 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_203
timestamp 0
transform 1 0 12374 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_54_207
timestamp 0
transform 1 0 12558 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_209
timestamp 0
transform 1 0 12650 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_211
timestamp 0
transform 1 0 12742 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_219
timestamp 0
transform 1 0 13110 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_54_223
timestamp 0
transform 1 0 13294 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_54_249
timestamp 0
transform 1 0 14490 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_54_261
timestamp 0
transform 1 0 15042 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_54_269
timestamp 0
transform 1 0 15410 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_271
timestamp 0
transform 1 0 15502 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_279
timestamp 0
transform 1 0 15870 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_54_283
timestamp 0
transform 1 0 16054 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_285
timestamp 0
transform 1 0 16146 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_310
timestamp 0
transform 1 0 17296 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_318
timestamp 0
transform 1 0 17664 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_326
timestamp 0
transform 1 0 18032 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_54_331
timestamp 0
transform 1 0 18262 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_339
timestamp 0
transform 1 0 18630 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_347
timestamp 0
transform 1 0 18998 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_355
timestamp 0
transform 1 0 19366 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_363
timestamp 0
transform 1 0 19734 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_371
timestamp 0
transform 1 0 20102 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_379
timestamp 0
transform 1 0 20470 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_54_387
timestamp 0
transform 1 0 20838 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_389
timestamp 0
transform 1 0 20930 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_54_391
timestamp 0
transform 1 0 21022 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_54_419
timestamp 0
transform 1 0 22310 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_427
timestamp 0
transform 1 0 22678 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_435
timestamp 0
transform 1 0 23046 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_443
timestamp 0
transform 1 0 23414 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_54_447
timestamp 0
transform 1 0 23598 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_449
timestamp 0
transform 1 0 23690 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_451
timestamp 0
transform 1 0 23782 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_459
timestamp 0
transform 1 0 24150 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_467
timestamp 0
transform 1 0 24518 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_475
timestamp 0
transform 1 0 24886 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_483
timestamp 0
transform 1 0 25254 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_491
timestamp 0
transform 1 0 25622 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_499
timestamp 0
transform 1 0 25990 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_54_507
timestamp 0
transform 1 0 26358 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_509
timestamp 0
transform 1 0 26450 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_511
timestamp 0
transform 1 0 26542 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_519
timestamp 0
transform 1 0 26910 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_527
timestamp 0
transform 1 0 27278 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_535
timestamp 0
transform 1 0 27646 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_543
timestamp 0
transform 1 0 28014 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_551
timestamp 0
transform 1 0 28382 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_54_559
timestamp 0
transform 1 0 28750 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_54_567
timestamp 0
transform 1 0 29118 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_569
timestamp 0
transform 1 0 29210 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_54_571
timestamp 0
transform 1 0 29302 0 1 17952
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_54_579
timestamp 0
transform 1 0 29670 0 1 17952
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_54_583
timestamp 0
transform 1 0 29854 0 1 17952
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_54_585
timestamp 0
transform 1 0 29946 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_55_0
timestamp 0
transform 1 0 3036 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_55_4
timestamp 0
transform 1 0 3220 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_55_30
timestamp 0
transform 1 0 4416 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_38
timestamp 0
transform 1 0 4784 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_46
timestamp 0
transform 1 0 5152 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_55_54
timestamp 0
transform 1 0 5520 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_55_58
timestamp 0
transform 1 0 5704 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_55_61
timestamp 0
transform 1 0 5842 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_55_74
timestamp 0
transform 1 0 6440 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_55_78
timestamp 0
transform 1 0 6624 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_55_103
timestamp 0
transform 1 0 7774 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_111
timestamp 0
transform 1 0 8142 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_55_119
timestamp 0
transform 1 0 8510 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_55_121
timestamp 0
transform 1 0 8602 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_129
timestamp 0
transform 1 0 8970 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_55_145
timestamp 0
transform 1 0 9706 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_55_149
timestamp 0
transform 1 0 9890 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_55_175
timestamp 0
transform 1 0 11086 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_55_179
timestamp 0
transform 1 0 11270 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_55_181
timestamp 0
transform 1 0 11362 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_189
timestamp 0
transform 1 0 11730 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_197
timestamp 0
transform 1 0 12098 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_55_205
timestamp 0
transform 1 0 12466 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_55_209
timestamp 0
transform 1 0 12650 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_55_211
timestamp 0
transform 1 0 12742 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_55_236
timestamp 0
transform 1 0 13892 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_55_241
timestamp 0
transform 1 0 14122 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_249
timestamp 0
transform 1 0 14490 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_55_257
timestamp 0
transform 1 0 14858 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_55_261
timestamp 0
transform 1 0 15042 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_55_263
timestamp 0
transform 1 0 15134 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_55_288
timestamp 0
transform 1 0 16284 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_55_295
timestamp 0
transform 1 0 16606 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_55_299
timestamp 0
transform 1 0 16790 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_55_301
timestamp 0
transform 1 0 16882 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_55_311
timestamp 0
transform 1 0 17342 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_319
timestamp 0
transform 1 0 17710 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_55_327
timestamp 0
transform 1 0 18078 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_55_331
timestamp 0
transform 1 0 18262 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_55_356
timestamp 0
transform 1 0 19412 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_55_361
timestamp 0
transform 1 0 19642 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_369
timestamp 0
transform 1 0 20010 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_377
timestamp 0
transform 1 0 20378 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_409
timestamp 0
transform 1 0 21850 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_55_417
timestamp 0
transform 1 0 22218 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_55_419
timestamp 0
transform 1 0 22310 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_55_421
timestamp 0
transform 1 0 22402 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_55_429
timestamp 0
transform 1 0 22770 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_55_433
timestamp 0
transform 1 0 22954 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_55_458
timestamp 0
transform 1 0 24104 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_55_468
timestamp 0
transform 1 0 24564 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_55_476
timestamp 0
transform 1 0 24932 0 -1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_55_481
timestamp 0
transform 1 0 25162 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_489
timestamp 0
transform 1 0 25530 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_497
timestamp 0
transform 1 0 25898 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_505
timestamp 0
transform 1 0 26266 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_513
timestamp 0
transform 1 0 26634 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_521
timestamp 0
transform 1 0 27002 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_55_529
timestamp 0
transform 1 0 27370 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_55_537
timestamp 0
transform 1 0 27738 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_55_539
timestamp 0
transform 1 0 27830 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_55_541
timestamp 0
transform 1 0 27922 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_55_549
timestamp 0
transform 1 0 28290 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_55_575
timestamp 0
transform 1 0 29486 0 -1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_55_583
timestamp 0
transform 1 0 29854 0 -1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_55_585
timestamp 0
transform 1 0 29946 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_56_0
timestamp 0
transform 1 0 3036 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_8
timestamp 0
transform 1 0 3404 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_16
timestamp 0
transform 1 0 3772 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_24
timestamp 0
transform 1 0 4140 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_28
timestamp 0
transform 1 0 4324 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_56_31
timestamp 0
transform 1 0 4462 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_56_41
timestamp 0
transform 1 0 4922 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_45
timestamp 0
transform 1 0 5106 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_56_47
timestamp 0
transform 1 0 5198 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_56_72
timestamp 0
transform 1 0 6348 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_80
timestamp 0
transform 1 0 6716 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_56_88
timestamp 0
transform 1 0 7084 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_56_91
timestamp 0
transform 1 0 7222 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_99
timestamp 0
transform 1 0 7590 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_107
timestamp 0
transform 1 0 7958 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_111
timestamp 0
transform 1 0 8142 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_56_113
timestamp 0
transform 1 0 8234 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_56_138
timestamp 0
transform 1 0 9384 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_146
timestamp 0
transform 1 0 9752 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_56_151
timestamp 0
transform 1 0 9982 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_159
timestamp 0
transform 1 0 10350 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_56_167
timestamp 0
transform 1 0 10718 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_56_169
timestamp 0
transform 1 0 10810 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_56_176
timestamp 0
transform 1 0 11132 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_180
timestamp 0
transform 1 0 11316 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_56_206
timestamp 0
transform 1 0 12512 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_56_211
timestamp 0
transform 1 0 12742 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_56_221
timestamp 0
transform 1 0 13202 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_229
timestamp 0
transform 1 0 13570 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_237
timestamp 0
transform 1 0 13938 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_56_241
timestamp 0
transform 1 0 14122 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_56_266
timestamp 0
transform 1 0 15272 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_56_271
timestamp 0
transform 1 0 15502 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_56_280
timestamp 0
transform 1 0 15916 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_56_284
timestamp 0
transform 1 0 16100 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_56_309
timestamp 0
transform 1 0 17250 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_317
timestamp 0
transform 1 0 17618 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_325
timestamp 0
transform 1 0 17986 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_56_329
timestamp 0
transform 1 0 18170 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_56_331
timestamp 0
transform 1 0 18262 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_339
timestamp 0
transform 1 0 18630 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_347
timestamp 0
transform 1 0 18998 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_56_351
timestamp 0
transform 1 0 19182 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_56_376
timestamp 0
transform 1 0 20332 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_56_386
timestamp 0
transform 1 0 20792 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_56_391
timestamp 0
transform 1 0 21022 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_56_400
timestamp 0
transform 1 0 21436 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_56_408
timestamp 0
transform 1 0 21804 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_56_410
timestamp 0
transform 1 0 21896 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_56_419
timestamp 0
transform 1 0 22310 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_427
timestamp 0
transform 1 0 22678 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_435
timestamp 0
transform 1 0 23046 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_443
timestamp 0
transform 1 0 23414 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_447
timestamp 0
transform 1 0 23598 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_56_449
timestamp 0
transform 1 0 23690 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_56_451
timestamp 0
transform 1 0 23782 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_56_459
timestamp 0
transform 1 0 24150 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_56_485
timestamp 0
transform 1 0 25346 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_493
timestamp 0
transform 1 0 25714 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_497
timestamp 0
transform 1 0 25898 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_56_506
timestamp 0
transform 1 0 26312 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_56_511
timestamp 0
transform 1 0 26542 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_56_519
timestamp 0
transform 1 0 26910 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_56_527
timestamp 0
transform 1 0 27278 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_56_535
timestamp 0
transform 1 0 27646 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_539
timestamp 0
transform 1 0 27830 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_56_541
timestamp 0
transform 1 0 27922 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_56_566
timestamp 0
transform 1 0 29072 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_56_571
timestamp 0
transform 1 0 29302 0 1 18496
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_56_579
timestamp 0
transform 1 0 29670 0 1 18496
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_56_583
timestamp 0
transform 1 0 29854 0 1 18496
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_56_585
timestamp 0
transform 1 0 29946 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_57_0
timestamp 0
transform 1 0 3036 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_57_32
timestamp 0
transform 1 0 4508 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_57_40
timestamp 0
transform 1 0 4876 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_48
timestamp 0
transform 1 0 5244 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_57_56
timestamp 0
transform 1 0 5612 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_57_61
timestamp 0
transform 1 0 5842 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 0
transform 1 0 6210 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_57_71
timestamp 0
transform 1 0 6302 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_57_79
timestamp 0
transform 1 0 6670 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_57_87
timestamp 0
transform 1 0 7038 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_57_91
timestamp 0
transform 1 0 7222 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_57_116
timestamp 0
transform 1 0 8372 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_57_121
timestamp 0
transform 1 0 8602 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_129
timestamp 0
transform 1 0 8970 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_137
timestamp 0
transform 1 0 9338 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_145
timestamp 0
transform 1 0 9706 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_153
timestamp 0
transform 1 0 10074 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_161
timestamp 0
transform 1 0 10442 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_169
timestamp 0
transform 1 0 10810 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_57_177
timestamp 0
transform 1 0 11178 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_57_179
timestamp 0
transform 1 0 11270 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_57_181
timestamp 0
transform 1 0 11362 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_57_189
timestamp 0
transform 1 0 11730 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_57_215
timestamp 0
transform 1 0 12926 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_223
timestamp 0
transform 1 0 13294 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_231
timestamp 0
transform 1 0 13662 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_57_239
timestamp 0
transform 1 0 14030 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_57_241
timestamp 0
transform 1 0 14122 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_57_269
timestamp 0
transform 1 0 15410 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_57_279
timestamp 0
transform 1 0 15870 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_287
timestamp 0
transform 1 0 16238 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_57_295
timestamp 0
transform 1 0 16606 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_57_299
timestamp 0
transform 1 0 16790 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_57_301
timestamp 0
transform 1 0 16882 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_309
timestamp 0
transform 1 0 17250 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_57_317
timestamp 0
transform 1 0 17618 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_57_342
timestamp 0
transform 1 0 18768 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_350
timestamp 0
transform 1 0 19136 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_57_358
timestamp 0
transform 1 0 19504 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_57_361
timestamp 0
transform 1 0 19642 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_369
timestamp 0
transform 1 0 20010 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_377
timestamp 0
transform 1 0 20378 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_385
timestamp 0
transform 1 0 20746 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_393
timestamp 0
transform 1 0 21114 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_401
timestamp 0
transform 1 0 21482 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_57_409
timestamp 0
transform 1 0 21850 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_57_417
timestamp 0
transform 1 0 22218 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_57_419
timestamp 0
transform 1 0 22310 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_57_421
timestamp 0
transform 1 0 22402 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_57_429
timestamp 0
transform 1 0 22770 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_57_431
timestamp 0
transform 1 0 22862 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_57_456
timestamp 0
transform 1 0 24012 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_57_467
timestamp 0
transform 1 0 24518 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_57_476
timestamp 0
transform 1 0 24932 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_57_481
timestamp 0
transform 1 0 25162 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_57_491
timestamp 0
transform 1 0 25622 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_57_499
timestamp 0
transform 1 0 25990 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_57_503
timestamp 0
transform 1 0 26174 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_57_529
timestamp 0
transform 1 0 27370 0 -1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_57_537
timestamp 0
transform 1 0 27738 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_57_539
timestamp 0
transform 1 0 27830 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_57_541
timestamp 0
transform 1 0 27922 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_57_545
timestamp 0
transform 1 0 28106 0 -1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_57_571
timestamp 0
transform 1 0 29302 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_57_581
timestamp 0
transform 1 0 29762 0 -1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_57_585
timestamp 0
transform 1 0 29946 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_58_0
timestamp 0
transform 1 0 3036 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_58_26
timestamp 0
transform 1 0 4232 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_58_31
timestamp 0
transform 1 0 4462 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_39
timestamp 0
transform 1 0 4830 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_47
timestamp 0
transform 1 0 5198 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_58_51
timestamp 0
transform 1 0 5382 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_58_53
timestamp 0
transform 1 0 5474 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_58_78
timestamp 0
transform 1 0 6624 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_58_86
timestamp 0
transform 1 0 6992 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_58_91
timestamp 0
transform 1 0 7222 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_58_119
timestamp 0
transform 1 0 8510 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_127
timestamp 0
transform 1 0 8878 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_135
timestamp 0
transform 1 0 9246 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_143
timestamp 0
transform 1 0 9614 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_58_147
timestamp 0
transform 1 0 9798 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_58_149
timestamp 0
transform 1 0 9890 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_58_151
timestamp 0
transform 1 0 9982 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_159
timestamp 0
transform 1 0 10350 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_167
timestamp 0
transform 1 0 10718 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_175
timestamp 0
transform 1 0 11086 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_183
timestamp 0
transform 1 0 11454 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_191
timestamp 0
transform 1 0 11822 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_199
timestamp 0
transform 1 0 12190 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_58_207
timestamp 0
transform 1 0 12558 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_58_209
timestamp 0
transform 1 0 12650 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_58_211
timestamp 0
transform 1 0 12742 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_219
timestamp 0
transform 1 0 13110 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_227
timestamp 0
transform 1 0 13478 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_235
timestamp 0
transform 1 0 13846 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_243
timestamp 0
transform 1 0 14214 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_251
timestamp 0
transform 1 0 14582 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_259
timestamp 0
transform 1 0 14950 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_58_267
timestamp 0
transform 1 0 15318 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_58_269
timestamp 0
transform 1 0 15410 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_58_271
timestamp 0
transform 1 0 15502 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_279
timestamp 0
transform 1 0 15870 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_287
timestamp 0
transform 1 0 16238 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_295
timestamp 0
transform 1 0 16606 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_303
timestamp 0
transform 1 0 16974 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_311
timestamp 0
transform 1 0 17342 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_319
timestamp 0
transform 1 0 17710 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_58_327
timestamp 0
transform 1 0 18078 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_58_329
timestamp 0
transform 1 0 18170 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_58_331
timestamp 0
transform 1 0 18262 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_339
timestamp 0
transform 1 0 18630 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_58_343
timestamp 0
transform 1 0 18814 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_58_369
timestamp 0
transform 1 0 20010 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_377
timestamp 0
transform 1 0 20378 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_385
timestamp 0
transform 1 0 20746 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_58_389
timestamp 0
transform 1 0 20930 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_58_391
timestamp 0
transform 1 0 21022 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_58_399
timestamp 0
transform 1 0 21390 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_58_424
timestamp 0
transform 1 0 22540 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_432
timestamp 0
transform 1 0 22908 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_440
timestamp 0
transform 1 0 23276 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_58_448
timestamp 0
transform 1 0 23644 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_58_451
timestamp 0
transform 1 0 23782 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_459
timestamp 0
transform 1 0 24150 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_58_463
timestamp 0
transform 1 0 24334 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_58_488
timestamp 0
transform 1 0 25484 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_496
timestamp 0
transform 1 0 25852 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_504
timestamp 0
transform 1 0 26220 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_58_508
timestamp 0
transform 1 0 26404 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_58_511
timestamp 0
transform 1 0 26542 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_519
timestamp 0
transform 1 0 26910 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_58_523
timestamp 0
transform 1 0 27094 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_58_530
timestamp 0
transform 1 0 27416 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_538
timestamp 0
transform 1 0 27784 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_546
timestamp 0
transform 1 0 28152 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_554
timestamp 0
transform 1 0 28520 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_562
timestamp 0
transform 1 0 28888 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_58_571
timestamp 0
transform 1 0 29302 0 1 19040
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_58_579
timestamp 0
transform 1 0 29670 0 1 19040
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_58_583
timestamp 0
transform 1 0 29854 0 1 19040
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_58_585
timestamp 0
transform 1 0 29946 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_0
timestamp 0
transform 1 0 3036 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_59_8
timestamp 0
transform 1 0 3404 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_10
timestamp 0
transform 1 0 3496 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_59_35
timestamp 0
transform 1 0 4646 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_59_47
timestamp 0
transform 1 0 5198 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_59_55
timestamp 0
transform 1 0 5566 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_59_59
timestamp 0
transform 1 0 5750 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_61
timestamp 0
transform 1 0 5842 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_69
timestamp 0
transform 1 0 6210 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_77
timestamp 0
transform 1 0 6578 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_59_85
timestamp 0
transform 1 0 6946 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_59_89
timestamp 0
transform 1 0 7130 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_91
timestamp 0
transform 1 0 7222 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_59_116
timestamp 0
transform 1 0 8372 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_59_121
timestamp 0
transform 1 0 8602 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_59_133
timestamp 0
transform 1 0 9154 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_141
timestamp 0
transform 1 0 9522 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_149
timestamp 0
transform 1 0 9890 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_157
timestamp 0
transform 1 0 10258 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_165
timestamp 0
transform 1 0 10626 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_59_173
timestamp 0
transform 1 0 10994 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_59_177
timestamp 0
transform 1 0 11178 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_179
timestamp 0
transform 1 0 11270 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_181
timestamp 0
transform 1 0 11362 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_189
timestamp 0
transform 1 0 11730 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_197
timestamp 0
transform 1 0 12098 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_205
timestamp 0
transform 1 0 12466 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_213
timestamp 0
transform 1 0 12834 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_221
timestamp 0
transform 1 0 13202 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_229
timestamp 0
transform 1 0 13570 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_59_237
timestamp 0
transform 1 0 13938 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_239
timestamp 0
transform 1 0 14030 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_241
timestamp 0
transform 1 0 14122 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_249
timestamp 0
transform 1 0 14490 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_257
timestamp 0
transform 1 0 14858 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_265
timestamp 0
transform 1 0 15226 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_273
timestamp 0
transform 1 0 15594 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_281
timestamp 0
transform 1 0 15962 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_289
timestamp 0
transform 1 0 16330 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_59_297
timestamp 0
transform 1 0 16698 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_299
timestamp 0
transform 1 0 16790 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_301
timestamp 0
transform 1 0 16882 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_309
timestamp 0
transform 1 0 17250 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_317
timestamp 0
transform 1 0 17618 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_325
timestamp 0
transform 1 0 17986 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_333
timestamp 0
transform 1 0 18354 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_341
timestamp 0
transform 1 0 18722 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_349
timestamp 0
transform 1 0 19090 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_59_357
timestamp 0
transform 1 0 19458 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_359
timestamp 0
transform 1 0 19550 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_361
timestamp 0
transform 1 0 19642 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_59_369
timestamp 0
transform 1 0 20010 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_59_373
timestamp 0
transform 1 0 20194 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_59_382
timestamp 0
transform 1 0 20608 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 0
transform 1 0 20976 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_59_416
timestamp 0
transform 1 0 22172 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_59_421
timestamp 0
transform 1 0 22402 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_59_433
timestamp 0
transform 1 0 22954 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_59_461
timestamp 0
transform 1 0 24242 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_469
timestamp 0
transform 1 0 24610 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_59_477
timestamp 0
transform 1 0 24978 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_479
timestamp 0
transform 1 0 25070 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_481
timestamp 0
transform 1 0 25162 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_489
timestamp 0
transform 1 0 25530 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_497
timestamp 0
transform 1 0 25898 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_505
timestamp 0
transform 1 0 26266 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_513
timestamp 0
transform 1 0 26634 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_521
timestamp 0
transform 1 0 27002 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_529
timestamp 0
transform 1 0 27370 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_59_537
timestamp 0
transform 1 0 27738 0 -1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_59_539
timestamp 0
transform 1 0 27830 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_59_541
timestamp 0
transform 1 0 27922 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_549
timestamp 0
transform 1 0 28290 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_557
timestamp 0
transform 1 0 28658 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_565
timestamp 0
transform 1 0 29026 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_59_573
timestamp 0
transform 1 0 29394 0 -1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_59_581
timestamp 0
transform 1 0 29762 0 -1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_59_585
timestamp 0
transform 1 0 29946 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_0
timestamp 0
transform 1 0 3036 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_8
timestamp 0
transform 1 0 3404 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_16
timestamp 0
transform 1 0 3772 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_24
timestamp 0
transform 1 0 4140 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_28
timestamp 0
transform 1 0 4324 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_60_31
timestamp 0
transform 1 0 4462 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_39
timestamp 0
transform 1 0 4830 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_47
timestamp 0
transform 1 0 5198 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_60_75
timestamp 0
transform 1 0 6486 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_83
timestamp 0
transform 1 0 6854 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_87
timestamp 0
transform 1 0 7038 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_60_89
timestamp 0
transform 1 0 7130 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_91
timestamp 0
transform 1 0 7222 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_99
timestamp 0
transform 1 0 7590 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_107
timestamp 0
transform 1 0 7958 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_115
timestamp 0
transform 1 0 8326 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_119
timestamp 0
transform 1 0 8510 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_60_121
timestamp 0
transform 1 0 8602 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_60_146
timestamp 0
transform 1 0 9752 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_60_151
timestamp 0
transform 1 0 9982 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_60_155
timestamp 0
transform 1 0 10166 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_60_165
timestamp 0
transform 1 0 10626 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_169
timestamp 0
transform 1 0 10810 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_60_171
timestamp 0
transform 1 0 10902 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_196
timestamp 0
transform 1 0 12052 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_204
timestamp 0
transform 1 0 12420 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_208
timestamp 0
transform 1 0 12604 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_60_211
timestamp 0
transform 1 0 12742 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_60_215
timestamp 0
transform 1 0 12926 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_240
timestamp 0
transform 1 0 14076 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_248
timestamp 0
transform 1 0 14444 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_256
timestamp 0
transform 1 0 14812 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_264
timestamp 0
transform 1 0 15180 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_268
timestamp 0
transform 1 0 15364 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_60_271
timestamp 0
transform 1 0 15502 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_60_279
timestamp 0
transform 1 0 15870 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_60_305
timestamp 0
transform 1 0 17066 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_313
timestamp 0
transform 1 0 17434 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_321
timestamp 0
transform 1 0 17802 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_60_329
timestamp 0
transform 1 0 18170 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_331
timestamp 0
transform 1 0 18262 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_339
timestamp 0
transform 1 0 18630 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_347
timestamp 0
transform 1 0 18998 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_379
timestamp 0
transform 1 0 20470 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_60_387
timestamp 0
transform 1 0 20838 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_60_389
timestamp 0
transform 1 0 20930 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_60_391
timestamp 0
transform 1 0 21022 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_395
timestamp 0
transform 1 0 21206 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_60_421
timestamp 0
transform 1 0 22402 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_429
timestamp 0
transform 1 0 22770 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_437
timestamp 0
transform 1 0 23138 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_445
timestamp 0
transform 1 0 23506 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_60_449
timestamp 0
transform 1 0 23690 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_451
timestamp 0
transform 1 0 23782 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_459
timestamp 0
transform 1 0 24150 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_467
timestamp 0
transform 1 0 24518 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_475
timestamp 0
transform 1 0 24886 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_483
timestamp 0
transform 1 0 25254 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_491
timestamp 0
transform 1 0 25622 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_499
timestamp 0
transform 1 0 25990 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_60_507
timestamp 0
transform 1 0 26358 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_60_509
timestamp 0
transform 1 0 26450 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_511
timestamp 0
transform 1 0 26542 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_519
timestamp 0
transform 1 0 26910 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_527
timestamp 0
transform 1 0 27278 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_535
timestamp 0
transform 1 0 27646 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_543
timestamp 0
transform 1 0 28014 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_551
timestamp 0
transform 1 0 28382 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_60_559
timestamp 0
transform 1 0 28750 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_60_567
timestamp 0
transform 1 0 29118 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_60_569
timestamp 0
transform 1 0 29210 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_60_571
timestamp 0
transform 1 0 29302 0 1 19584
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_60_579
timestamp 0
transform 1 0 29670 0 1 19584
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_60_583
timestamp 0
transform 1 0 29854 0 1 19584
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_60_585
timestamp 0
transform 1 0 29946 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_61_0
timestamp 0
transform 1 0 3036 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_8
timestamp 0
transform 1 0 3404 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_16
timestamp 0
transform 1 0 3772 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_24
timestamp 0
transform 1 0 4140 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_32
timestamp 0
transform 1 0 4508 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_40
timestamp 0
transform 1 0 4876 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_48
timestamp 0
transform 1 0 5244 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_56
timestamp 0
transform 1 0 5612 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_61_61
timestamp 0
transform 1 0 5842 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_61_65
timestamp 0
transform 1 0 6026 0 -1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_61_67
timestamp 0
transform 1 0 6118 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_61_92
timestamp 0
transform 1 0 7268 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_100
timestamp 0
transform 1 0 7636 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_108
timestamp 0
transform 1 0 8004 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_116
timestamp 0
transform 1 0 8372 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_61_121
timestamp 0
transform 1 0 8602 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_61_149
timestamp 0
transform 1 0 9890 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_61_159
timestamp 0
transform 1 0 10350 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_167
timestamp 0
transform 1 0 10718 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_175
timestamp 0
transform 1 0 11086 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_61_179
timestamp 0
transform 1 0 11270 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_61_181
timestamp 0
transform 1 0 11362 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_196
timestamp 0
transform 1 0 12052 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_61_207
timestamp 0
transform 1 0 12558 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_61_211
timestamp 0
transform 1 0 12742 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_61_236
timestamp 0
transform 1 0 13892 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_61_241
timestamp 0
transform 1 0 14122 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_249
timestamp 0
transform 1 0 14490 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_257
timestamp 0
transform 1 0 14858 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_265
timestamp 0
transform 1 0 15226 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_61_269
timestamp 0
transform 1 0 15410 0 -1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_61_271
timestamp 0
transform 1 0 15502 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_61_296
timestamp 0
transform 1 0 16652 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_61_301
timestamp 0
transform 1 0 16882 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_309
timestamp 0
transform 1 0 17250 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_61_317
timestamp 0
transform 1 0 17618 0 -1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_61_343
timestamp 0
transform 1 0 18814 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_61_350
timestamp 0
transform 1 0 19136 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_61_358
timestamp 0
transform 1 0 19504 0 -1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_61_361
timestamp 0
transform 1 0 19642 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_369
timestamp 0
transform 1 0 20010 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_377
timestamp 0
transform 1 0 20378 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_61_381
timestamp 0
transform 1 0 20562 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_61_389
timestamp 0
transform 1 0 20930 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_397
timestamp 0
transform 1 0 21298 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_405
timestamp 0
transform 1 0 21666 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_413
timestamp 0
transform 1 0 22034 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_61_417
timestamp 0
transform 1 0 22218 0 -1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_61_419
timestamp 0
transform 1 0 22310 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_61_421
timestamp 0
transform 1 0 22402 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_429
timestamp 0
transform 1 0 22770 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_61_433
timestamp 0
transform 1 0 22954 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_61_458
timestamp 0
transform 1 0 24104 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_61_468
timestamp 0
transform 1 0 24564 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_476
timestamp 0
transform 1 0 24932 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_61_481
timestamp 0
transform 1 0 25162 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_61_489
timestamp 0
transform 1 0 25530 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_61_514
timestamp 0
transform 1 0 26680 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_522
timestamp 0
transform 1 0 27048 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_530
timestamp 0
transform 1 0 27416 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_61_538
timestamp 0
transform 1 0 27784 0 -1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_61_541
timestamp 0
transform 1 0 27922 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_549
timestamp 0
transform 1 0 28290 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_557
timestamp 0
transform 1 0 28658 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_565
timestamp 0
transform 1 0 29026 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_61_573
timestamp 0
transform 1 0 29394 0 -1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_61_581
timestamp 0
transform 1 0 29762 0 -1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_61_585
timestamp 0
transform 1 0 29946 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_62_0
timestamp 0
transform 1 0 3036 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_8
timestamp 0
transform 1 0 3404 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_16
timestamp 0
transform 1 0 3772 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_62_24
timestamp 0
transform 1 0 4140 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_62_28
timestamp 0
transform 1 0 4324 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_62_31
timestamp 0
transform 1 0 4462 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_39
timestamp 0
transform 1 0 4830 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_47
timestamp 0
transform 1 0 5198 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_49
timestamp 0
transform 1 0 5290 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_62_74
timestamp 0
transform 1 0 6440 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_82
timestamp 0
transform 1 0 6808 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_91
timestamp 0
transform 1 0 7222 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_99
timestamp 0
transform 1 0 7590 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_107
timestamp 0
transform 1 0 7958 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_115
timestamp 0
transform 1 0 8326 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_123
timestamp 0
transform 1 0 8694 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_131
timestamp 0
transform 1 0 9062 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_139
timestamp 0
transform 1 0 9430 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_147
timestamp 0
transform 1 0 9798 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_149
timestamp 0
transform 1 0 9890 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_62_151
timestamp 0
transform 1 0 9982 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_159
timestamp 0
transform 1 0 10350 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_167
timestamp 0
transform 1 0 10718 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_62_175
timestamp 0
transform 1 0 11086 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_62_179
timestamp 0
transform 1 0 11270 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_181
timestamp 0
transform 1 0 11362 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_62_206
timestamp 0
transform 1 0 12512 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_62_211
timestamp 0
transform 1 0 12742 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_62_239
timestamp 0
transform 1 0 14030 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_62_251
timestamp 0
transform 1 0 14582 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_259
timestamp 0
transform 1 0 14950 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_267
timestamp 0
transform 1 0 15318 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_269
timestamp 0
transform 1 0 15410 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_62_271
timestamp 0
transform 1 0 15502 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_279
timestamp 0
transform 1 0 15870 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_62_305
timestamp 0
transform 1 0 17066 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_62_317
timestamp 0
transform 1 0 17618 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_62_325
timestamp 0
transform 1 0 17986 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_62_329
timestamp 0
transform 1 0 18170 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_62_331
timestamp 0
transform 1 0 18262 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_339
timestamp 0
transform 1 0 18630 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_347
timestamp 0
transform 1 0 18998 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_355
timestamp 0
transform 1 0 19366 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_357
timestamp 0
transform 1 0 19458 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_62_382
timestamp 0
transform 1 0 20608 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_391
timestamp 0
transform 1 0 21022 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_399
timestamp 0
transform 1 0 21390 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_407
timestamp 0
transform 1 0 21758 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_415
timestamp 0
transform 1 0 22126 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_423
timestamp 0
transform 1 0 22494 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_431
timestamp 0
transform 1 0 22862 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_439
timestamp 0
transform 1 0 23230 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_447
timestamp 0
transform 1 0 23598 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_449
timestamp 0
transform 1 0 23690 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_62_451
timestamp 0
transform 1 0 23782 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_459
timestamp 0
transform 1 0 24150 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_467
timestamp 0
transform 1 0 24518 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_475
timestamp 0
transform 1 0 24886 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_483
timestamp 0
transform 1 0 25254 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_491
timestamp 0
transform 1 0 25622 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_499
timestamp 0
transform 1 0 25990 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_507
timestamp 0
transform 1 0 26358 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_509
timestamp 0
transform 1 0 26450 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_62_511
timestamp 0
transform 1 0 26542 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_62_523
timestamp 0
transform 1 0 27094 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_62_531
timestamp 0
transform 1 0 27462 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_62_539
timestamp 0
transform 1 0 27830 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_541
timestamp 0
transform 1 0 27922 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_62_566
timestamp 0
transform 1 0 29072 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_62_571
timestamp 0
transform 1 0 29302 0 1 20128
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_62_579
timestamp 0
transform 1 0 29670 0 1 20128
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_62_583
timestamp 0
transform 1 0 29854 0 1 20128
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_62_585
timestamp 0
transform 1 0 29946 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_63_0
timestamp 0
transform 1 0 3036 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_8
timestamp 0
transform 1 0 3404 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_40
timestamp 0
transform 1 0 4876 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_48
timestamp 0
transform 1 0 5244 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_56
timestamp 0
transform 1 0 5612 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_63_61
timestamp 0
transform 1 0 5842 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_63_69
timestamp 0
transform 1 0 6210 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_63_71
timestamp 0
transform 1 0 6302 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_63_96
timestamp 0
transform 1 0 7452 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_63_107
timestamp 0
transform 1 0 7958 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_115
timestamp 0
transform 1 0 8326 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_63_119
timestamp 0
transform 1 0 8510 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_63_121
timestamp 0
transform 1 0 8602 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_129
timestamp 0
transform 1 0 8970 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_137
timestamp 0
transform 1 0 9338 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_145
timestamp 0
transform 1 0 9706 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_153
timestamp 0
transform 1 0 10074 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_161
timestamp 0
transform 1 0 10442 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_169
timestamp 0
transform 1 0 10810 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_63_177
timestamp 0
transform 1 0 11178 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_63_179
timestamp 0
transform 1 0 11270 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_63_181
timestamp 0
transform 1 0 11362 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_63_209
timestamp 0
transform 1 0 12650 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_217
timestamp 0
transform 1 0 13018 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_225
timestamp 0
transform 1 0 13386 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_233
timestamp 0
transform 1 0 13754 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_63_237
timestamp 0
transform 1 0 13938 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_63_239
timestamp 0
transform 1 0 14030 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_63_241
timestamp 0
transform 1 0 14122 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_249
timestamp 0
transform 1 0 14490 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_63_253
timestamp 0
transform 1 0 14674 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_63_258
timestamp 0
transform 1 0 14904 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_63_262
timestamp 0
transform 1 0 15088 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_63_264
timestamp 0
transform 1 0 15180 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_63_272
timestamp 0
transform 1 0 15548 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_280
timestamp 0
transform 1 0 15916 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_288
timestamp 0
transform 1 0 16284 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_296
timestamp 0
transform 1 0 16652 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_63_301
timestamp 0
transform 1 0 16882 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_309
timestamp 0
transform 1 0 17250 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_317
timestamp 0
transform 1 0 17618 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_325
timestamp 0
transform 1 0 17986 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_333
timestamp 0
transform 1 0 18354 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_341
timestamp 0
transform 1 0 18722 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_349
timestamp 0
transform 1 0 19090 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_63_357
timestamp 0
transform 1 0 19458 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_63_359
timestamp 0
transform 1 0 19550 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_63_361
timestamp 0
transform 1 0 19642 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_369
timestamp 0
transform 1 0 20010 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_377
timestamp 0
transform 1 0 20378 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_385
timestamp 0
transform 1 0 20746 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_63_389
timestamp 0
transform 1 0 20930 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 0
transform 1 0 21022 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_63_416
timestamp 0
transform 1 0 22172 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_63_421
timestamp 0
transform 1 0 22402 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_63_431
timestamp 0
transform 1 0 22862 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_439
timestamp 0
transform 1 0 23230 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_63_443
timestamp 0
transform 1 0 23414 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_63_469
timestamp 0
transform 1 0 24610 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_63_477
timestamp 0
transform 1 0 24978 0 -1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_63_479
timestamp 0
transform 1 0 25070 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_63_481
timestamp 0
transform 1 0 25162 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_513
timestamp 0
transform 1 0 26634 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_63_520
timestamp 0
transform 1 0 26956 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_63_528
timestamp 0
transform 1 0 27324 0 -1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_63_536
timestamp 0
transform 1 0 27692 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_63_541
timestamp 0
transform 1 0 27922 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_63_569
timestamp 0
transform 1 0 29210 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_63_581
timestamp 0
transform 1 0 29762 0 -1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_63_585
timestamp 0
transform 1 0 29946 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_64_0
timestamp 0
transform 1 0 3036 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_64_26
timestamp 0
transform 1 0 4232 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_64_31
timestamp 0
transform 1 0 4462 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_39
timestamp 0
transform 1 0 4830 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_64_47
timestamp 0
transform 1 0 5198 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_64_51
timestamp 0
transform 1 0 5382 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_64_53
timestamp 0
transform 1 0 5474 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_64_78
timestamp 0
transform 1 0 6624 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_64_86
timestamp 0
transform 1 0 6992 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_64_91
timestamp 0
transform 1 0 7222 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_123
timestamp 0
transform 1 0 8694 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_131
timestamp 0
transform 1 0 9062 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_139
timestamp 0
transform 1 0 9430 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_64_147
timestamp 0
transform 1 0 9798 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 0
transform 1 0 9890 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_64_151
timestamp 0
transform 1 0 9982 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_159
timestamp 0
transform 1 0 10350 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_64_167
timestamp 0
transform 1 0 10718 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_64_193
timestamp 0
transform 1 0 11914 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_201
timestamp 0
transform 1 0 12282 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_64_209
timestamp 0
transform 1 0 12650 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_64_211
timestamp 0
transform 1 0 12742 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_219
timestamp 0
transform 1 0 13110 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_251
timestamp 0
transform 1 0 14582 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_259
timestamp 0
transform 1 0 14950 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_64_267
timestamp 0
transform 1 0 15318 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_64_269
timestamp 0
transform 1 0 15410 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_64_271
timestamp 0
transform 1 0 15502 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_279
timestamp 0
transform 1 0 15870 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_287
timestamp 0
transform 1 0 16238 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_295
timestamp 0
transform 1 0 16606 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_303
timestamp 0
transform 1 0 16974 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_311
timestamp 0
transform 1 0 17342 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_319
timestamp 0
transform 1 0 17710 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_64_327
timestamp 0
transform 1 0 18078 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_64_329
timestamp 0
transform 1 0 18170 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_64_331
timestamp 0
transform 1 0 18262 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_339
timestamp 0
transform 1 0 18630 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_371
timestamp 0
transform 1 0 20102 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_379
timestamp 0
transform 1 0 20470 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_64_387
timestamp 0
transform 1 0 20838 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_64_389
timestamp 0
transform 1 0 20930 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_64_391
timestamp 0
transform 1 0 21022 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_64_419
timestamp 0
transform 1 0 22310 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_64_432
timestamp 0
transform 1 0 22908 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_440
timestamp 0
transform 1 0 23276 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_64_448
timestamp 0
transform 1 0 23644 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_64_451
timestamp 0
transform 1 0 23782 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_459
timestamp 0
transform 1 0 24150 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_64_467
timestamp 0
transform 1 0 24518 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_64_474
timestamp 0
transform 1 0 24840 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_482
timestamp 0
transform 1 0 25208 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_490
timestamp 0
transform 1 0 25576 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_498
timestamp 0
transform 1 0 25944 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_64_506
timestamp 0
transform 1 0 26312 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_64_511
timestamp 0
transform 1 0 26542 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_519
timestamp 0
transform 1 0 26910 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_64_527
timestamp 0
transform 1 0 27278 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_64_535
timestamp 0
transform 1 0 27646 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_64_539
timestamp 0
transform 1 0 27830 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_64_541
timestamp 0
transform 1 0 27922 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_64_566
timestamp 0
transform 1 0 29072 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_64_571
timestamp 0
transform 1 0 29302 0 1 20672
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_64_579
timestamp 0
transform 1 0 29670 0 1 20672
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_64_583
timestamp 0
transform 1 0 29854 0 1 20672
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_64_585
timestamp 0
transform 1 0 29946 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_65_0
timestamp 0
transform 1 0 3036 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_65_8
timestamp 0
transform 1 0 3404 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_65_34
timestamp 0
transform 1 0 4600 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_65_44
timestamp 0
transform 1 0 5060 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_52
timestamp 0
transform 1 0 5428 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_61
timestamp 0
transform 1 0 5842 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_69
timestamp 0
transform 1 0 6210 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_65_73
timestamp 0
transform 1 0 6394 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_65_82
timestamp 0
transform 1 0 6808 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_65_90
timestamp 0
transform 1 0 7176 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_65_116
timestamp 0
transform 1 0 8372 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_65_121
timestamp 0
transform 1 0 8602 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_129
timestamp 0
transform 1 0 8970 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_137
timestamp 0
transform 1 0 9338 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_65_165
timestamp 0
transform 1 0 10626 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_173
timestamp 0
transform 1 0 10994 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_65_177
timestamp 0
transform 1 0 11178 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_65_179
timestamp 0
transform 1 0 11270 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_65_181
timestamp 0
transform 1 0 11362 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_189
timestamp 0
transform 1 0 11730 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_197
timestamp 0
transform 1 0 12098 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_65_201
timestamp 0
transform 1 0 12282 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_65_211
timestamp 0
transform 1 0 12742 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_219
timestamp 0
transform 1 0 13110 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_227
timestamp 0
transform 1 0 13478 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_235
timestamp 0
transform 1 0 13846 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_65_239
timestamp 0
transform 1 0 14030 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_65_241
timestamp 0
transform 1 0 14122 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_249
timestamp 0
transform 1 0 14490 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_257
timestamp 0
transform 1 0 14858 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_265
timestamp 0
transform 1 0 15226 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_273
timestamp 0
transform 1 0 15594 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_281
timestamp 0
transform 1 0 15962 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_289
timestamp 0
transform 1 0 16330 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_65_297
timestamp 0
transform 1 0 16698 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_65_299
timestamp 0
transform 1 0 16790 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_65_301
timestamp 0
transform 1 0 16882 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_309
timestamp 0
transform 1 0 17250 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_317
timestamp 0
transform 1 0 17618 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_325
timestamp 0
transform 1 0 17986 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_65_329
timestamp 0
transform 1 0 18170 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_65_331
timestamp 0
transform 1 0 18262 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_65_356
timestamp 0
transform 1 0 19412 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_65_361
timestamp 0
transform 1 0 19642 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_65_369
timestamp 0
transform 1 0 20010 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_65_379
timestamp 0
transform 1 0 20470 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_387
timestamp 0
transform 1 0 20838 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_395
timestamp 0
transform 1 0 21206 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_403
timestamp 0
transform 1 0 21574 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_411
timestamp 0
transform 1 0 21942 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_65_419
timestamp 0
transform 1 0 22310 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_65_421
timestamp 0
transform 1 0 22402 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_429
timestamp 0
transform 1 0 22770 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_437
timestamp 0
transform 1 0 23138 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_65_441
timestamp 0
transform 1 0 23322 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_65_467
timestamp 0
transform 1 0 24518 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_475
timestamp 0
transform 1 0 24886 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_65_479
timestamp 0
transform 1 0 25070 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_65_481
timestamp 0
transform 1 0 25162 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_489
timestamp 0
transform 1 0 25530 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_65_493
timestamp 0
transform 1 0 25714 0 -1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_65_519
timestamp 0
transform 1 0 26910 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_527
timestamp 0
transform 1 0 27278 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_535
timestamp 0
transform 1 0 27646 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_65_539
timestamp 0
transform 1 0 27830 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_65_541
timestamp 0
transform 1 0 27922 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_549
timestamp 0
transform 1 0 28290 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_557
timestamp 0
transform 1 0 28658 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_565
timestamp 0
transform 1 0 29026 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_65_573
timestamp 0
transform 1 0 29394 0 -1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_65_581
timestamp 0
transform 1 0 29762 0 -1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_65_585
timestamp 0
transform 1 0 29946 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_0
timestamp 0
transform 1 0 3036 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_8
timestamp 0
transform 1 0 3404 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_16
timestamp 0
transform 1 0 3772 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_66_24
timestamp 0
transform 1 0 4140 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_66_28
timestamp 0
transform 1 0 4324 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_66_31
timestamp 0
transform 1 0 4462 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_66_41
timestamp 0
transform 1 0 4922 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_73
timestamp 0
transform 1 0 6394 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_81
timestamp 0
transform 1 0 6762 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_66_89
timestamp 0
transform 1 0 7130 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_91
timestamp 0
transform 1 0 7222 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_99
timestamp 0
transform 1 0 7590 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_66_107
timestamp 0
transform 1 0 7958 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_109
timestamp 0
transform 1 0 8050 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_66_118
timestamp 0
transform 1 0 8464 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_66_146
timestamp 0
transform 1 0 9752 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_66_151
timestamp 0
transform 1 0 9982 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_66_159
timestamp 0
transform 1 0 10350 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_66_163
timestamp 0
transform 1 0 10534 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_171
timestamp 0
transform 1 0 10902 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_66_179
timestamp 0
transform 1 0 11270 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_181
timestamp 0
transform 1 0 11362 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_66_206
timestamp 0
transform 1 0 12512 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_66_211
timestamp 0
transform 1 0 12742 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_219
timestamp 0
transform 1 0 13110 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_227
timestamp 0
transform 1 0 13478 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_66_235
timestamp 0
transform 1 0 13846 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_66_239
timestamp 0
transform 1 0 14030 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_241
timestamp 0
transform 1 0 14122 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_66_266
timestamp 0
transform 1 0 15272 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_66_271
timestamp 0
transform 1 0 15502 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_279
timestamp 0
transform 1 0 15870 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_66_287
timestamp 0
transform 1 0 16238 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_289
timestamp 0
transform 1 0 16330 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_301
timestamp 0
transform 1 0 16882 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_309
timestamp 0
transform 1 0 17250 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_317
timestamp 0
transform 1 0 17618 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_66_325
timestamp 0
transform 1 0 17986 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_66_329
timestamp 0
transform 1 0 18170 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_331
timestamp 0
transform 1 0 18262 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_339
timestamp 0
transform 1 0 18630 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_66_347
timestamp 0
transform 1 0 18998 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_66_351
timestamp 0
transform 1 0 19182 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_353
timestamp 0
transform 1 0 19274 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_378
timestamp 0
transform 1 0 20424 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_66_386
timestamp 0
transform 1 0 20792 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_66_391
timestamp 0
transform 1 0 21022 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_399
timestamp 0
transform 1 0 21390 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_407
timestamp 0
transform 1 0 21758 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_415
timestamp 0
transform 1 0 22126 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_423
timestamp 0
transform 1 0 22494 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_431
timestamp 0
transform 1 0 22862 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_439
timestamp 0
transform 1 0 23230 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_66_447
timestamp 0
transform 1 0 23598 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_449
timestamp 0
transform 1 0 23690 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_451
timestamp 0
transform 1 0 23782 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_459
timestamp 0
transform 1 0 24150 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_467
timestamp 0
transform 1 0 24518 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_475
timestamp 0
transform 1 0 24886 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_483
timestamp 0
transform 1 0 25254 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_491
timestamp 0
transform 1 0 25622 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_499
timestamp 0
transform 1 0 25990 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_66_507
timestamp 0
transform 1 0 26358 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_509
timestamp 0
transform 1 0 26450 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_511
timestamp 0
transform 1 0 26542 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_519
timestamp 0
transform 1 0 26910 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_527
timestamp 0
transform 1 0 27278 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_535
timestamp 0
transform 1 0 27646 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_543
timestamp 0
transform 1 0 28014 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_551
timestamp 0
transform 1 0 28382 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_66_559
timestamp 0
transform 1 0 28750 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_66_567
timestamp 0
transform 1 0 29118 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_569
timestamp 0
transform 1 0 29210 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_66_571
timestamp 0
transform 1 0 29302 0 1 21216
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_66_579
timestamp 0
transform 1 0 29670 0 1 21216
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_66_583
timestamp 0
transform 1 0 29854 0 1 21216
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_66_585
timestamp 0
transform 1 0 29946 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_0
timestamp 0
transform 1 0 3036 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_32
timestamp 0
transform 1 0 4508 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_67_36
timestamp 0
transform 1 0 4692 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_41
timestamp 0
transform 1 0 4922 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_49
timestamp 0
transform 1 0 5290 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 0
transform 1 0 5658 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_67_59
timestamp 0
transform 1 0 5750 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_61
timestamp 0
transform 1 0 5842 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_69
timestamp 0
transform 1 0 6210 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_67_81
timestamp 0
transform 1 0 6762 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_67_89
timestamp 0
transform 1 0 7130 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_67_91
timestamp 0
transform 1 0 7222 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_67_116
timestamp 0
transform 1 0 8372 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_67_121
timestamp 0
transform 1 0 8602 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_129
timestamp 0
transform 1 0 8970 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_137
timestamp 0
transform 1 0 9338 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_67_141
timestamp 0
transform 1 0 9522 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_67_143
timestamp 0
transform 1 0 9614 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_168
timestamp 0
transform 1 0 10764 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_176
timestamp 0
transform 1 0 11132 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_67_181
timestamp 0
transform 1 0 11362 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_67_185
timestamp 0
transform 1 0 11546 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_67_211
timestamp 0
transform 1 0 12742 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_67_224
timestamp 0
transform 1 0 13340 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_232
timestamp 0
transform 1 0 13708 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_241
timestamp 0
transform 1 0 14122 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_67_269
timestamp 0
transform 1 0 15410 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_67_290
timestamp 0
transform 1 0 16376 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_67_298
timestamp 0
transform 1 0 16744 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_67_301
timestamp 0
transform 1 0 16882 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_309
timestamp 0
transform 1 0 17250 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_67_313
timestamp 0
transform 1 0 17434 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_67_325
timestamp 0
transform 1 0 17986 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_67_337
timestamp 0
transform 1 0 18538 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_345
timestamp 0
transform 1 0 18906 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_353
timestamp 0
transform 1 0 19274 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_67_357
timestamp 0
transform 1 0 19458 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_67_359
timestamp 0
transform 1 0 19550 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_361
timestamp 0
transform 1 0 19642 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_369
timestamp 0
transform 1 0 20010 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_377
timestamp 0
transform 1 0 20378 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_385
timestamp 0
transform 1 0 20746 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_393
timestamp 0
transform 1 0 21114 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_401
timestamp 0
transform 1 0 21482 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_409
timestamp 0
transform 1 0 21850 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_67_417
timestamp 0
transform 1 0 22218 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_67_419
timestamp 0
transform 1 0 22310 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_421
timestamp 0
transform 1 0 22402 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_429
timestamp 0
transform 1 0 22770 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_437
timestamp 0
transform 1 0 23138 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_445
timestamp 0
transform 1 0 23506 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_453
timestamp 0
transform 1 0 23874 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_461
timestamp 0
transform 1 0 24242 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_469
timestamp 0
transform 1 0 24610 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_67_477
timestamp 0
transform 1 0 24978 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_67_479
timestamp 0
transform 1 0 25070 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_481
timestamp 0
transform 1 0 25162 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_67_489
timestamp 0
transform 1 0 25530 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_497
timestamp 0
transform 1 0 25898 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_67_501
timestamp 0
transform 1 0 26082 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_67_526
timestamp 0
transform 1 0 27232 0 -1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_67_534
timestamp 0
transform 1 0 27600 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_67_538
timestamp 0
transform 1 0 27784 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_67_541
timestamp 0
transform 1 0 27922 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_67_545
timestamp 0
transform 1 0 28106 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_67_571
timestamp 0
transform 1 0 29302 0 -1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_67_583
timestamp 0
transform 1 0 29854 0 -1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_67_585
timestamp 0
transform 1 0 29946 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_68_0
timestamp 0
transform 1 0 3036 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_8
timestamp 0
transform 1 0 3404 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_16
timestamp 0
transform 1 0 3772 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_68_24
timestamp 0
transform 1 0 4140 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_68_28
timestamp 0
transform 1 0 4324 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_68_31
timestamp 0
transform 1 0 4462 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_68_39
timestamp 0
transform 1 0 4830 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_68_43
timestamp 0
transform 1 0 5014 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_68_45
timestamp 0
transform 1 0 5106 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_68_70
timestamp 0
transform 1 0 6256 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_68_81
timestamp 0
transform 1 0 6762 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_68_89
timestamp 0
transform 1 0 7130 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_68_91
timestamp 0
transform 1 0 7222 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_99
timestamp 0
transform 1 0 7590 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_107
timestamp 0
transform 1 0 7958 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_115
timestamp 0
transform 1 0 8326 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_123
timestamp 0
transform 1 0 8694 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_131
timestamp 0
transform 1 0 9062 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_139
timestamp 0
transform 1 0 9430 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_68_147
timestamp 0
transform 1 0 9798 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_68_149
timestamp 0
transform 1 0 9890 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_68_151
timestamp 0
transform 1 0 9982 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_68_162
timestamp 0
transform 1 0 10488 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_170
timestamp 0
transform 1 0 10856 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_68_178
timestamp 0
transform 1 0 11224 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_68_204
timestamp 0
transform 1 0 12420 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_68_208
timestamp 0
transform 1 0 12604 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_68_211
timestamp 0
transform 1 0 12742 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_219
timestamp 0
transform 1 0 13110 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_227
timestamp 0
transform 1 0 13478 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_235
timestamp 0
transform 1 0 13846 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_68_243
timestamp 0
transform 1 0 14214 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_68_253
timestamp 0
transform 1 0 14674 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_68_266
timestamp 0
transform 1 0 15272 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_68_271
timestamp 0
transform 1 0 15502 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_279
timestamp 0
transform 1 0 15870 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_68_287
timestamp 0
transform 1 0 16238 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_68_296
timestamp 0
transform 1 0 16652 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_68_308
timestamp 0
transform 1 0 17204 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_68_312
timestamp 0
transform 1 0 17388 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_68_314
timestamp 0
transform 1 0 17480 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_68_326
timestamp 0
transform 1 0 18032 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_68_331
timestamp 0
transform 1 0 18262 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_339
timestamp 0
transform 1 0 18630 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_347
timestamp 0
transform 1 0 18998 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_68_355
timestamp 0
transform 1 0 19366 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_68_357
timestamp 0
transform 1 0 19458 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_68_382
timestamp 0
transform 1 0 20608 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_68_391
timestamp 0
transform 1 0 21022 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_68_419
timestamp 0
transform 1 0 22310 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_68_431
timestamp 0
transform 1 0 22862 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_442
timestamp 0
transform 1 0 23368 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_451
timestamp 0
transform 1 0 23782 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_68_459
timestamp 0
transform 1 0 24150 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_68_463
timestamp 0
transform 1 0 24334 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_68_489
timestamp 0
transform 1 0 25530 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_68_497
timestamp 0
transform 1 0 25898 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_68_505
timestamp 0
transform 1 0 26266 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_68_509
timestamp 0
transform 1 0 26450 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_68_511
timestamp 0
transform 1 0 26542 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_68_539
timestamp 0
transform 1 0 27830 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_68_551
timestamp 0
transform 1 0 28382 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_68_559
timestamp 0
transform 1 0 28750 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_68_567
timestamp 0
transform 1 0 29118 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_68_569
timestamp 0
transform 1 0 29210 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_68_571
timestamp 0
transform 1 0 29302 0 1 21760
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_68_579
timestamp 0
transform 1 0 29670 0 1 21760
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_68_583
timestamp 0
transform 1 0 29854 0 1 21760
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_68_585
timestamp 0
transform 1 0 29946 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_0
timestamp 0
transform 1 0 3036 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_69_8
timestamp 0
transform 1 0 3404 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_69_34
timestamp 0
transform 1 0 4600 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_42
timestamp 0
transform 1 0 4968 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_50
timestamp 0
transform 1 0 5336 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_69_58
timestamp 0
transform 1 0 5704 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_69_61
timestamp 0
transform 1 0 5842 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_69
timestamp 0
transform 1 0 6210 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_77
timestamp 0
transform 1 0 6578 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_69_85
timestamp 0
transform 1 0 6946 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_69_89
timestamp 0
transform 1 0 7130 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_69_115
timestamp 0
transform 1 0 8326 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_69_119
timestamp 0
transform 1 0 8510 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_121
timestamp 0
transform 1 0 8602 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_69_129
timestamp 0
transform 1 0 8970 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_69_131
timestamp 0
transform 1 0 9062 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_156
timestamp 0
transform 1 0 10212 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_164
timestamp 0
transform 1 0 10580 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_172
timestamp 0
transform 1 0 10948 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_181
timestamp 0
transform 1 0 11362 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_189
timestamp 0
transform 1 0 11730 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_197
timestamp 0
transform 1 0 12098 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_205
timestamp 0
transform 1 0 12466 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_213
timestamp 0
transform 1 0 12834 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_221
timestamp 0
transform 1 0 13202 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_229
timestamp 0
transform 1 0 13570 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_69_237
timestamp 0
transform 1 0 13938 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_69_239
timestamp 0
transform 1 0 14030 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_241
timestamp 0
transform 1 0 14122 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_249
timestamp 0
transform 1 0 14490 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_69_257
timestamp 0
transform 1 0 14858 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_267
timestamp 0
transform 1 0 15318 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_275
timestamp 0
transform 1 0 15686 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_69_283
timestamp 0
transform 1 0 16054 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_69_293
timestamp 0
transform 1 0 16514 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_69_297
timestamp 0
transform 1 0 16698 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_69_299
timestamp 0
transform 1 0 16790 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_301
timestamp 0
transform 1 0 16882 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_309
timestamp 0
transform 1 0 17250 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_328
timestamp 0
transform 1 0 18124 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_340
timestamp 0
transform 1 0 18676 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_348
timestamp 0
transform 1 0 19044 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_69_356
timestamp 0
transform 1 0 19412 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_69_361
timestamp 0
transform 1 0 19642 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_369
timestamp 0
transform 1 0 20010 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_377
timestamp 0
transform 1 0 20378 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_69_385
timestamp 0
transform 1 0 20746 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_69_389
timestamp 0
transform 1 0 20930 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 0
transform 1 0 21022 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_69_416
timestamp 0
transform 1 0 22172 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_69_421
timestamp 0
transform 1 0 22402 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_429
timestamp 0
transform 1 0 22770 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_69_437
timestamp 0
transform 1 0 23138 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_69_439
timestamp 0
transform 1 0 23230 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_69_456
timestamp 0
transform 1 0 24012 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_69_464
timestamp 0
transform 1 0 24380 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_69_472
timestamp 0
transform 1 0 24748 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_69_481
timestamp 0
transform 1 0 25162 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_69_485
timestamp 0
transform 1 0 25346 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_493
timestamp 0
transform 1 0 25714 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_69_501
timestamp 0
transform 1 0 26082 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_69_527
timestamp 0
transform 1 0 27278 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_69_535
timestamp 0
transform 1 0 27646 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_69_539
timestamp 0
transform 1 0 27830 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_69_541
timestamp 0
transform 1 0 27922 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_69_545
timestamp 0
transform 1 0 28106 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_69_547
timestamp 0
transform 1 0 28198 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_69_572
timestamp 0
transform 1 0 29348 0 -1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_69_580
timestamp 0
transform 1 0 29716 0 -1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_69_584
timestamp 0
transform 1 0 29900 0 -1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_2  FILLER_70_0
timestamp 0
transform 1 0 3036 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_70_26
timestamp 0
transform 1 0 4232 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_70_31
timestamp 0
transform 1 0 4462 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_70_43
timestamp 0
transform 1 0 5014 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_47
timestamp 0
transform 1 0 5198 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_70_73
timestamp 0
transform 1 0 6394 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_81
timestamp 0
transform 1 0 6762 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_70_89
timestamp 0
transform 1 0 7130 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_70_91
timestamp 0
transform 1 0 7222 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_70_119
timestamp 0
transform 1 0 8510 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_70_131
timestamp 0
transform 1 0 9062 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_139
timestamp 0
transform 1 0 9430 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_70_147
timestamp 0
transform 1 0 9798 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_70_149
timestamp 0
transform 1 0 9890 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_70_151
timestamp 0
transform 1 0 9982 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_159
timestamp 0
transform 1 0 10350 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_167
timestamp 0
transform 1 0 10718 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_175
timestamp 0
transform 1 0 11086 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_183
timestamp 0
transform 1 0 11454 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_191
timestamp 0
transform 1 0 11822 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_199
timestamp 0
transform 1 0 12190 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_70_207
timestamp 0
transform 1 0 12558 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_70_209
timestamp 0
transform 1 0 12650 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_70_211
timestamp 0
transform 1 0 12742 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_219
timestamp 0
transform 1 0 13110 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_223
timestamp 0
transform 1 0 13294 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_70_234
timestamp 0
transform 1 0 13800 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_242
timestamp 0
transform 1 0 14168 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_250
timestamp 0
transform 1 0 14536 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_70_254
timestamp 0
transform 1 0 14720 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_70_264
timestamp 0
transform 1 0 15180 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_268
timestamp 0
transform 1 0 15364 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_70_271
timestamp 0
transform 1 0 15502 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_279
timestamp 0
transform 1 0 15870 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_283
timestamp 0
transform 1 0 16054 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_70_294
timestamp 0
transform 1 0 16560 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_302
timestamp 0
transform 1 0 16928 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_310
timestamp 0
transform 1 0 17296 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_314
timestamp 0
transform 1 0 17480 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_70_316
timestamp 0
transform 1 0 17572 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_70_322
timestamp 0
transform 1 0 17848 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_331
timestamp 0
transform 1 0 18262 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_70_351
timestamp 0
transform 1 0 19182 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_359
timestamp 0
transform 1 0 19550 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_367
timestamp 0
transform 1 0 19918 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_375
timestamp 0
transform 1 0 20286 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_383
timestamp 0
transform 1 0 20654 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_387
timestamp 0
transform 1 0 20838 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_70_389
timestamp 0
transform 1 0 20930 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_70_391
timestamp 0
transform 1 0 21022 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_395
timestamp 0
transform 1 0 21206 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_70_421
timestamp 0
transform 1 0 22402 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_429
timestamp 0
transform 1 0 22770 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_70_436
timestamp 0
transform 1 0 23092 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_70_443
timestamp 0
transform 1 0 23414 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_447
timestamp 0
transform 1 0 23598 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_70_449
timestamp 0
transform 1 0 23690 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_70_451
timestamp 0
transform 1 0 23782 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_459
timestamp 0
transform 1 0 24150 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_70_463
timestamp 0
transform 1 0 24334 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_70_488
timestamp 0
transform 1 0 25484 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_496
timestamp 0
transform 1 0 25852 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_504
timestamp 0
transform 1 0 26220 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_508
timestamp 0
transform 1 0 26404 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_70_511
timestamp 0
transform 1 0 26542 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_519
timestamp 0
transform 1 0 26910 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_527
timestamp 0
transform 1 0 27278 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_535
timestamp 0
transform 1 0 27646 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_543
timestamp 0
transform 1 0 28014 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_551
timestamp 0
transform 1 0 28382 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_70_559
timestamp 0
transform 1 0 28750 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_70_567
timestamp 0
transform 1 0 29118 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_70_569
timestamp 0
transform 1 0 29210 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_70_571
timestamp 0
transform 1 0 29302 0 1 22304
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_70_579
timestamp 0
transform 1 0 29670 0 1 22304
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_70_583
timestamp 0
transform 1 0 29854 0 1 22304
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_70_585
timestamp 0
transform 1 0 29946 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_71_0
timestamp 0
transform 1 0 3036 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_32
timestamp 0
transform 1 0 4508 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_40
timestamp 0
transform 1 0 4876 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_48
timestamp 0
transform 1 0 5244 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_56
timestamp 0
transform 1 0 5612 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_71_61
timestamp 0
transform 1 0 5842 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_69
timestamp 0
transform 1 0 6210 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_77
timestamp 0
transform 1 0 6578 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_85
timestamp 0
transform 1 0 6946 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_89
timestamp 0
transform 1 0 7130 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_91
timestamp 0
transform 1 0 7222 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_71_116
timestamp 0
transform 1 0 8372 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_71_121
timestamp 0
transform 1 0 8602 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_129
timestamp 0
transform 1 0 8970 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_137
timestamp 0
transform 1 0 9338 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_145
timestamp 0
transform 1 0 9706 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_149
timestamp 0
transform 1 0 9890 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_151
timestamp 0
transform 1 0 9982 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_71_176
timestamp 0
transform 1 0 11132 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_71_181
timestamp 0
transform 1 0 11362 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_189
timestamp 0
transform 1 0 11730 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_197
timestamp 0
transform 1 0 12098 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_205
timestamp 0
transform 1 0 12466 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_209
timestamp 0
transform 1 0 12650 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_211
timestamp 0
transform 1 0 12742 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_71_221
timestamp 0
transform 1 0 13202 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_71_234
timestamp 0
transform 1 0 13800 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_238
timestamp 0
transform 1 0 13984 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_71_241
timestamp 0
transform 1 0 14122 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_71_249
timestamp 0
transform 1 0 14490 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_251
timestamp 0
transform 1 0 14582 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_71_261
timestamp 0
transform 1 0 15042 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_269
timestamp 0
transform 1 0 15410 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_273
timestamp 0
transform 1 0 15594 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_275
timestamp 0
transform 1 0 15686 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_71_285
timestamp 0
transform 1 0 16146 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_293
timestamp 0
transform 1 0 16514 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_297
timestamp 0
transform 1 0 16698 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_299
timestamp 0
transform 1 0 16790 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_71_301
timestamp 0
transform 1 0 16882 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_309
timestamp 0
transform 1 0 17250 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_333
timestamp 0
transform 1 0 18354 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_71_341
timestamp 0
transform 1 0 18722 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_356
timestamp 0
transform 1 0 19412 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_71_361
timestamp 0
transform 1 0 19642 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_365
timestamp 0
transform 1 0 19826 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_367
timestamp 0
transform 1 0 19918 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_71_375
timestamp 0
transform 1 0 20286 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_383
timestamp 0
transform 1 0 20654 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_391
timestamp 0
transform 1 0 21022 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_399
timestamp 0
transform 1 0 21390 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_407
timestamp 0
transform 1 0 21758 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_415
timestamp 0
transform 1 0 22126 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_71_419
timestamp 0
transform 1 0 22310 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_71_421
timestamp 0
transform 1 0 22402 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_429
timestamp 0
transform 1 0 22770 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_71_437
timestamp 0
transform 1 0 23138 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_71_455
timestamp 0
transform 1 0 23966 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_71_463
timestamp 0
transform 1 0 24334 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_471
timestamp 0
transform 1 0 24702 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_71_479
timestamp 0
transform 1 0 25070 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_71_481
timestamp 0
transform 1 0 25162 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_489
timestamp 0
transform 1 0 25530 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_497
timestamp 0
transform 1 0 25898 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_505
timestamp 0
transform 1 0 26266 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_513
timestamp 0
transform 1 0 26634 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_521
timestamp 0
transform 1 0 27002 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_71_529
timestamp 0
transform 1 0 27370 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_71_537
timestamp 0
transform 1 0 27738 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_539
timestamp 0
transform 1 0 27830 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_71_541
timestamp 0
transform 1 0 27922 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_545
timestamp 0
transform 1 0 28106 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_71_571
timestamp 0
transform 1 0 29302 0 -1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_71_579
timestamp 0
transform 1 0 29670 0 -1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_71_583
timestamp 0
transform 1 0 29854 0 -1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_71_585
timestamp 0
transform 1 0 29946 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_0
timestamp 0
transform 1 0 3036 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_8
timestamp 0
transform 1 0 3404 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_16
timestamp 0
transform 1 0 3772 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_24
timestamp 0
transform 1 0 4140 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_72_28
timestamp 0
transform 1 0 4324 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_72_31
timestamp 0
transform 1 0 4462 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_39
timestamp 0
transform 1 0 4830 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_47
timestamp 0
transform 1 0 5198 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_72_51
timestamp 0
transform 1 0 5382 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_72_77
timestamp 0
transform 1 0 6578 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_85
timestamp 0
transform 1 0 6946 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_72_89
timestamp 0
transform 1 0 7130 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_91
timestamp 0
transform 1 0 7222 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_99
timestamp 0
transform 1 0 7590 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_107
timestamp 0
transform 1 0 7958 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_115
timestamp 0
transform 1 0 8326 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_123
timestamp 0
transform 1 0 8694 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_131
timestamp 0
transform 1 0 9062 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_72_135
timestamp 0
transform 1 0 9246 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_139
timestamp 0
transform 1 0 9430 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_72_147
timestamp 0
transform 1 0 9798 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_72_149
timestamp 0
transform 1 0 9890 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_151
timestamp 0
transform 1 0 9982 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_159
timestamp 0
transform 1 0 10350 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_167
timestamp 0
transform 1 0 10718 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_199
timestamp 0
transform 1 0 12190 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_72_207
timestamp 0
transform 1 0 12558 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_72_209
timestamp 0
transform 1 0 12650 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_211
timestamp 0
transform 1 0 12742 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_219
timestamp 0
transform 1 0 13110 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_72_223
timestamp 0
transform 1 0 13294 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_233
timestamp 0
transform 1 0 13754 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_241
timestamp 0
transform 1 0 14122 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_249
timestamp 0
transform 1 0 14490 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 0
transform 1 0 14674 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_72_255
timestamp 0
transform 1 0 14766 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_72_265
timestamp 0
transform 1 0 15226 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_72_269
timestamp 0
transform 1 0 15410 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_271
timestamp 0
transform 1 0 15502 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_72_279
timestamp 0
transform 1 0 15870 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_72_290
timestamp 0
transform 1 0 16376 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_72_294
timestamp 0
transform 1 0 16560 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_304
timestamp 0
transform 1 0 17020 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_72_312
timestamp 0
transform 1 0 17388 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_72_317
timestamp 0
transform 1 0 17618 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_72_325
timestamp 0
transform 1 0 17986 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_72_329
timestamp 0
transform 1 0 18170 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_331
timestamp 0
transform 1 0 18262 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_339
timestamp 0
transform 1 0 18630 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_347
timestamp 0
transform 1 0 18998 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_355
timestamp 0
transform 1 0 19366 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_72_359
timestamp 0
transform 1 0 19550 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_72_367
timestamp 0
transform 1 0 19918 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_72_384
timestamp 0
transform 1 0 20700 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_72_388
timestamp 0
transform 1 0 20884 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_72_391
timestamp 0
transform 1 0 21022 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_72_399
timestamp 0
transform 1 0 21390 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_72_407
timestamp 0
transform 1 0 21758 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_415
timestamp 0
transform 1 0 22126 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_72_419
timestamp 0
transform 1 0 22310 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_72_421
timestamp 0
transform 1 0 22402 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_72_429
timestamp 0
transform 1 0 22770 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_72_436
timestamp 0
transform 1 0 23092 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_444
timestamp 0
transform 1 0 23460 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_72_448
timestamp 0
transform 1 0 23644 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_72_451
timestamp 0
transform 1 0 23782 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_459
timestamp 0
transform 1 0 24150 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_72_467
timestamp 0
transform 1 0 24518 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_72_493
timestamp 0
transform 1 0 25714 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_501
timestamp 0
transform 1 0 26082 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_72_509
timestamp 0
transform 1 0 26450 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_511
timestamp 0
transform 1 0 26542 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_519
timestamp 0
transform 1 0 26910 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_527
timestamp 0
transform 1 0 27278 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_535
timestamp 0
transform 1 0 27646 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_543
timestamp 0
transform 1 0 28014 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_551
timestamp 0
transform 1 0 28382 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_72_559
timestamp 0
transform 1 0 28750 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_72_567
timestamp 0
transform 1 0 29118 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_72_569
timestamp 0
transform 1 0 29210 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_72_571
timestamp 0
transform 1 0 29302 0 1 22848
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_72_579
timestamp 0
transform 1 0 29670 0 1 22848
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_72_583
timestamp 0
transform 1 0 29854 0 1 22848
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_72_585
timestamp 0
transform 1 0 29946 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_0
timestamp 0
transform 1 0 3036 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_8
timestamp 0
transform 1 0 3404 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_16
timestamp 0
transform 1 0 3772 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_24
timestamp 0
transform 1 0 4140 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_32
timestamp 0
transform 1 0 4508 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_40
timestamp 0
transform 1 0 4876 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_48
timestamp 0
transform 1 0 5244 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_73_56
timestamp 0
transform 1 0 5612 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_73_61
timestamp 0
transform 1 0 5842 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_73_69
timestamp 0
transform 1 0 6210 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_76
timestamp 0
transform 1 0 6532 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_84
timestamp 0
transform 1 0 6900 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_92
timestamp 0
transform 1 0 7268 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_100
timestamp 0
transform 1 0 7636 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_108
timestamp 0
transform 1 0 8004 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_73_116
timestamp 0
transform 1 0 8372 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_73_121
timestamp 0
transform 1 0 8602 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_73_129
timestamp 0
transform 1 0 8970 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_73_133
timestamp 0
transform 1 0 9154 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_73_158
timestamp 0
transform 1 0 10304 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_73_162
timestamp 0
transform 1 0 10488 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_164
timestamp 0
transform 1 0 10580 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_170
timestamp 0
transform 1 0 10856 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_73_178
timestamp 0
transform 1 0 11224 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_73_181
timestamp 0
transform 1 0 11362 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_73_188
timestamp 0
transform 1 0 11684 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_73_192
timestamp 0
transform 1 0 11868 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_194
timestamp 0
transform 1 0 11960 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_201
timestamp 0
transform 1 0 12282 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_73_209
timestamp 0
transform 1 0 12650 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_73_213
timestamp 0
transform 1 0 12834 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_215
timestamp 0
transform 1 0 12926 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_225
timestamp 0
transform 1 0 13386 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_73_233
timestamp 0
transform 1 0 13754 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_73_237
timestamp 0
transform 1 0 13938 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_239
timestamp 0
transform 1 0 14030 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_241
timestamp 0
transform 1 0 14122 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_73_249
timestamp 0
transform 1 0 14490 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_73_260
timestamp 0
transform 1 0 14996 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_268
timestamp 0
transform 1 0 15364 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_276
timestamp 0
transform 1 0 15732 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_73_284
timestamp 0
transform 1 0 16100 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_286
timestamp 0
transform 1 0 16192 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_73_296
timestamp 0
transform 1 0 16652 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_73_301
timestamp 0
transform 1 0 16882 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_73_313
timestamp 0
transform 1 0 17434 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_73_321
timestamp 0
transform 1 0 17802 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_73_332
timestamp 0
transform 1 0 18308 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_73_340
timestamp 0
transform 1 0 18676 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_73_344
timestamp 0
transform 1 0 18860 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_346
timestamp 0
transform 1 0 18952 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_73_356
timestamp 0
transform 1 0 19412 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_73_361
timestamp 0
transform 1 0 19642 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_369
timestamp 0
transform 1 0 20010 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_73_377
timestamp 0
transform 1 0 20378 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_73_394
timestamp 0
transform 1 0 21160 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_73_414
timestamp 0
transform 1 0 22080 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_73_418
timestamp 0
transform 1 0 22264 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_73_421
timestamp 0
transform 1 0 22402 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_429
timestamp 0
transform 1 0 22770 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_437
timestamp 0
transform 1 0 23138 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_445
timestamp 0
transform 1 0 23506 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_453
timestamp 0
transform 1 0 23874 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_461
timestamp 0
transform 1 0 24242 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_469
timestamp 0
transform 1 0 24610 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_73_477
timestamp 0
transform 1 0 24978 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_479
timestamp 0
transform 1 0 25070 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_481
timestamp 0
transform 1 0 25162 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_489
timestamp 0
transform 1 0 25530 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_497
timestamp 0
transform 1 0 25898 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_505
timestamp 0
transform 1 0 26266 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_513
timestamp 0
transform 1 0 26634 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_521
timestamp 0
transform 1 0 27002 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_529
timestamp 0
transform 1 0 27370 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_73_537
timestamp 0
transform 1 0 27738 0 -1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_73_539
timestamp 0
transform 1 0 27830 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_73_541
timestamp 0
transform 1 0 27922 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_549
timestamp 0
transform 1 0 28290 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_557
timestamp 0
transform 1 0 28658 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_565
timestamp 0
transform 1 0 29026 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_73_573
timestamp 0
transform 1 0 29394 0 -1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_73_581
timestamp 0
transform 1 0 29762 0 -1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_73_585
timestamp 0
transform 1 0 29946 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_74_0
timestamp 0
transform 1 0 3036 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_8
timestamp 0
transform 1 0 3404 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_16
timestamp 0
transform 1 0 3772 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_24
timestamp 0
transform 1 0 4140 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_74_28
timestamp 0
transform 1 0 4324 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_74_31
timestamp 0
transform 1 0 4462 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_39
timestamp 0
transform 1 0 4830 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_74_43
timestamp 0
transform 1 0 5014 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_74_69
timestamp 0
transform 1 0 6210 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_74_80
timestamp 0
transform 1 0 6716 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_74_88
timestamp 0
transform 1 0 7084 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_74_91
timestamp 0
transform 1 0 7222 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_99
timestamp 0
transform 1 0 7590 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_107
timestamp 0
transform 1 0 7958 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_74_135
timestamp 0
transform 1 0 9246 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_74_142
timestamp 0
transform 1 0 9568 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_151
timestamp 0
transform 1 0 9982 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_74_162
timestamp 0
transform 1 0 10488 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_74_170
timestamp 0
transform 1 0 10856 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_74_172
timestamp 0
transform 1 0 10948 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_74_197
timestamp 0
transform 1 0 12098 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_205
timestamp 0
transform 1 0 12466 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_74_209
timestamp 0
transform 1 0 12650 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_74_211
timestamp 0
transform 1 0 12742 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_74_215
timestamp 0
transform 1 0 12926 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_74_225
timestamp 0
transform 1 0 13386 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_233
timestamp 0
transform 1 0 13754 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_241
timestamp 0
transform 1 0 14122 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_249
timestamp 0
transform 1 0 14490 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_257
timestamp 0
transform 1 0 14858 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_265
timestamp 0
transform 1 0 15226 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_74_269
timestamp 0
transform 1 0 15410 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_74_271
timestamp 0
transform 1 0 15502 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_279
timestamp 0
transform 1 0 15870 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_287
timestamp 0
transform 1 0 16238 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_295
timestamp 0
transform 1 0 16606 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_303
timestamp 0
transform 1 0 16974 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_311
timestamp 0
transform 1 0 17342 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_74_315
timestamp 0
transform 1 0 17526 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_74_317
timestamp 0
transform 1 0 17618 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_74_326
timestamp 0
transform 1 0 18032 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_74_331
timestamp 0
transform 1 0 18262 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_74_339
timestamp 0
transform 1 0 18630 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_347
timestamp 0
transform 1 0 18998 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_379
timestamp 0
transform 1 0 20470 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_74_387
timestamp 0
transform 1 0 20838 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_74_389
timestamp 0
transform 1 0 20930 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_74_391
timestamp 0
transform 1 0 21022 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_74_399
timestamp 0
transform 1 0 21390 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_74_407
timestamp 0
transform 1 0 21758 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_74_432
timestamp 0
transform 1 0 22908 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_74_443
timestamp 0
transform 1 0 23414 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_74_447
timestamp 0
transform 1 0 23598 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_74_449
timestamp 0
transform 1 0 23690 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_74_451
timestamp 0
transform 1 0 23782 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_74_459
timestamp 0
transform 1 0 24150 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_74_461
timestamp 0
transform 1 0 24242 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_74_478
timestamp 0
transform 1 0 25024 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_486
timestamp 0
transform 1 0 25392 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_494
timestamp 0
transform 1 0 25760 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_502
timestamp 0
transform 1 0 26128 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_511
timestamp 0
transform 1 0 26542 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_519
timestamp 0
transform 1 0 26910 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_527
timestamp 0
transform 1 0 27278 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_535
timestamp 0
transform 1 0 27646 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_543
timestamp 0
transform 1 0 28014 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_551
timestamp 0
transform 1 0 28382 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_74_559
timestamp 0
transform 1 0 28750 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_74_567
timestamp 0
transform 1 0 29118 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_74_569
timestamp 0
transform 1 0 29210 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_74_571
timestamp 0
transform 1 0 29302 0 1 23392
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_74_579
timestamp 0
transform 1 0 29670 0 1 23392
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_74_583
timestamp 0
transform 1 0 29854 0 1 23392
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_74_585
timestamp 0
transform 1 0 29946 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_0
timestamp 0
transform 1 0 3036 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_75_8
timestamp 0
transform 1 0 3404 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_75_33
timestamp 0
transform 1 0 4554 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_75_45
timestamp 0
transform 1 0 5106 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_75_53
timestamp 0
transform 1 0 5474 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_75_57
timestamp 0
transform 1 0 5658 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_75_59
timestamp 0
transform 1 0 5750 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_61
timestamp 0
transform 1 0 5842 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_75_69
timestamp 0
transform 1 0 6210 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_75_71
timestamp 0
transform 1 0 6302 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_76
timestamp 0
transform 1 0 6532 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_108
timestamp 0
transform 1 0 8004 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_75_116
timestamp 0
transform 1 0 8372 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_75_121
timestamp 0
transform 1 0 8602 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_75_129
timestamp 0
transform 1 0 8970 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_154
timestamp 0
transform 1 0 10120 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_162
timestamp 0
transform 1 0 10488 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_170
timestamp 0
transform 1 0 10856 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_75_178
timestamp 0
transform 1 0 11224 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_75_181
timestamp 0
transform 1 0 11362 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_189
timestamp 0
transform 1 0 11730 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_197
timestamp 0
transform 1 0 12098 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_205
timestamp 0
transform 1 0 12466 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_222
timestamp 0
transform 1 0 13248 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_230
timestamp 0
transform 1 0 13616 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_75_238
timestamp 0
transform 1 0 13984 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_75_241
timestamp 0
transform 1 0 14122 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_75_249
timestamp 0
transform 1 0 14490 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_75_253
timestamp 0
transform 1 0 14674 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_75_255
timestamp 0
transform 1 0 14766 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_265
timestamp 0
transform 1 0 15226 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_273
timestamp 0
transform 1 0 15594 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_281
timestamp 0
transform 1 0 15962 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_289
timestamp 0
transform 1 0 16330 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_75_297
timestamp 0
transform 1 0 16698 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_75_299
timestamp 0
transform 1 0 16790 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_301
timestamp 0
transform 1 0 16882 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_309
timestamp 0
transform 1 0 17250 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_75_317
timestamp 0
transform 1 0 17618 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_75_328
timestamp 0
transform 1 0 18124 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_75_348
timestamp 0
transform 1 0 19044 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_75_356
timestamp 0
transform 1 0 19412 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_75_361
timestamp 0
transform 1 0 19642 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_369
timestamp 0
transform 1 0 20010 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_377
timestamp 0
transform 1 0 20378 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_385
timestamp 0
transform 1 0 20746 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_75_393
timestamp 0
transform 1 0 21114 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_75_401
timestamp 0
transform 1 0 21482 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_409
timestamp 0
transform 1 0 21850 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_75_417
timestamp 0
transform 1 0 22218 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_75_419
timestamp 0
transform 1 0 22310 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_421
timestamp 0
transform 1 0 22402 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_429
timestamp 0
transform 1 0 22770 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_437
timestamp 0
transform 1 0 23138 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_75_445
timestamp 0
transform 1 0 23506 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_75_451
timestamp 0
transform 1 0 23782 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_75_471
timestamp 0
transform 1 0 24702 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_75_479
timestamp 0
transform 1 0 25070 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_481
timestamp 0
transform 1 0 25162 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_489
timestamp 0
transform 1 0 25530 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_497
timestamp 0
transform 1 0 25898 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_505
timestamp 0
transform 1 0 26266 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_513
timestamp 0
transform 1 0 26634 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_521
timestamp 0
transform 1 0 27002 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_529
timestamp 0
transform 1 0 27370 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_75_537
timestamp 0
transform 1 0 27738 0 -1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_75_539
timestamp 0
transform 1 0 27830 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_75_541
timestamp 0
transform 1 0 27922 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_549
timestamp 0
transform 1 0 28290 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_557
timestamp 0
transform 1 0 28658 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_565
timestamp 0
transform 1 0 29026 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_75_573
timestamp 0
transform 1 0 29394 0 -1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_75_581
timestamp 0
transform 1 0 29762 0 -1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_75_585
timestamp 0
transform 1 0 29946 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_76_0
timestamp 0
transform 1 0 3036 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_76_26
timestamp 0
transform 1 0 4232 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_76_31
timestamp 0
transform 1 0 4462 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_76_39
timestamp 0
transform 1 0 4830 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_76_41
timestamp 0
transform 1 0 4922 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_76_46
timestamp 0
transform 1 0 5152 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_54
timestamp 0
transform 1 0 5520 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_62
timestamp 0
transform 1 0 5888 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_70
timestamp 0
transform 1 0 6256 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_78
timestamp 0
transform 1 0 6624 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_86
timestamp 0
transform 1 0 6992 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_76_91
timestamp 0
transform 1 0 7222 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_99
timestamp 0
transform 1 0 7590 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_76_107
timestamp 0
transform 1 0 7958 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_76_133
timestamp 0
transform 1 0 9154 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_141
timestamp 0
transform 1 0 9522 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_76_149
timestamp 0
transform 1 0 9890 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_76_151
timestamp 0
transform 1 0 9982 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_159
timestamp 0
transform 1 0 10350 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_167
timestamp 0
transform 1 0 10718 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_175
timestamp 0
transform 1 0 11086 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_183
timestamp 0
transform 1 0 11454 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_191
timestamp 0
transform 1 0 11822 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_195
timestamp 0
transform 1 0 12006 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_76_197
timestamp 0
transform 1 0 12098 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_76_206
timestamp 0
transform 1 0 12512 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_76_211
timestamp 0
transform 1 0 12742 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_219
timestamp 0
transform 1 0 13110 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_227
timestamp 0
transform 1 0 13478 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_248
timestamp 0
transform 1 0 14444 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_256
timestamp 0
transform 1 0 14812 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_264
timestamp 0
transform 1 0 15180 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_268
timestamp 0
transform 1 0 15364 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_76_271
timestamp 0
transform 1 0 15502 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_279
timestamp 0
transform 1 0 15870 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_76_287
timestamp 0
transform 1 0 16238 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_76_294
timestamp 0
transform 1 0 16560 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_298
timestamp 0
transform 1 0 16744 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_76_308
timestamp 0
transform 1 0 17204 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_316
timestamp 0
transform 1 0 17572 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_324
timestamp 0
transform 1 0 17940 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_328
timestamp 0
transform 1 0 18124 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_76_331
timestamp 0
transform 1 0 18262 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_76_339
timestamp 0
transform 1 0 18630 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_347
timestamp 0
transform 1 0 18998 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_355
timestamp 0
transform 1 0 19366 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_363
timestamp 0
transform 1 0 19734 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_371
timestamp 0
transform 1 0 20102 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_375
timestamp 0
transform 1 0 20286 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_76_384
timestamp 0
transform 1 0 20700 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_388
timestamp 0
transform 1 0 20884 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_76_391
timestamp 0
transform 1 0 21022 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_399
timestamp 0
transform 1 0 21390 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_403
timestamp 0
transform 1 0 21574 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_76_405
timestamp 0
transform 1 0 21666 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_76_430
timestamp 0
transform 1 0 22816 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_438
timestamp 0
transform 1 0 23184 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_446
timestamp 0
transform 1 0 23552 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_76_451
timestamp 0
transform 1 0 23782 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_455
timestamp 0
transform 1 0 23966 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_76_457
timestamp 0
transform 1 0 24058 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_76_462
timestamp 0
transform 1 0 24288 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_76_470
timestamp 0
transform 1 0 24656 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_478
timestamp 0
transform 1 0 25024 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_486
timestamp 0
transform 1 0 25392 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_494
timestamp 0
transform 1 0 25760 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_502
timestamp 0
transform 1 0 26128 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_511
timestamp 0
transform 1 0 26542 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_519
timestamp 0
transform 1 0 26910 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_527
timestamp 0
transform 1 0 27278 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_535
timestamp 0
transform 1 0 27646 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_543
timestamp 0
transform 1 0 28014 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_551
timestamp 0
transform 1 0 28382 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_76_559
timestamp 0
transform 1 0 28750 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_76_567
timestamp 0
transform 1 0 29118 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_76_569
timestamp 0
transform 1 0 29210 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_76_571
timestamp 0
transform 1 0 29302 0 1 23936
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_76_579
timestamp 0
transform 1 0 29670 0 1 23936
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_76_583
timestamp 0
transform 1 0 29854 0 1 23936
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_76_585
timestamp 0
transform 1 0 29946 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_0
timestamp 0
transform 1 0 3036 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_77_8
timestamp 0
transform 1 0 3404 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_33
timestamp 0
transform 1 0 4554 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_41
timestamp 0
transform 1 0 4922 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_49
timestamp 0
transform 1 0 5290 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 0
transform 1 0 5658 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_59
timestamp 0
transform 1 0 5750 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_61
timestamp 0
transform 1 0 5842 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_69
timestamp 0
transform 1 0 6210 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_77
timestamp 0
transform 1 0 6578 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_77_81
timestamp 0
transform 1 0 6762 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_83
timestamp 0
transform 1 0 6854 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_108
timestamp 0
transform 1 0 8004 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_116
timestamp 0
transform 1 0 8372 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_77_121
timestamp 0
transform 1 0 8602 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_129
timestamp 0
transform 1 0 8970 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_77_139
timestamp 0
transform 1 0 9430 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_147
timestamp 0
transform 1 0 9798 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_155
timestamp 0
transform 1 0 10166 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_163
timestamp 0
transform 1 0 10534 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_171
timestamp 0
transform 1 0 10902 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_77_179
timestamp 0
transform 1 0 11270 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_181
timestamp 0
transform 1 0 11362 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_189
timestamp 0
transform 1 0 11730 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_77_193
timestamp 0
transform 1 0 11914 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_77_203
timestamp 0
transform 1 0 12374 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_211
timestamp 0
transform 1 0 12742 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_219
timestamp 0
transform 1 0 13110 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_227
timestamp 0
transform 1 0 13478 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_235
timestamp 0
transform 1 0 13846 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_77_239
timestamp 0
transform 1 0 14030 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_241
timestamp 0
transform 1 0 14122 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_249
timestamp 0
transform 1 0 14490 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_257
timestamp 0
transform 1 0 14858 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_265
timestamp 0
transform 1 0 15226 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_273
timestamp 0
transform 1 0 15594 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_77_277
timestamp 0
transform 1 0 15778 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 0
transform 1 0 15870 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_77_293
timestamp 0
transform 1 0 16514 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_77_297
timestamp 0
transform 1 0 16698 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_299
timestamp 0
transform 1 0 16790 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_301
timestamp 0
transform 1 0 16882 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_309
timestamp 0
transform 1 0 17250 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_77_313
timestamp 0
transform 1 0 17434 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_321
timestamp 0
transform 1 0 17802 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_329
timestamp 0
transform 1 0 18170 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_337
timestamp 0
transform 1 0 18538 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_345
timestamp 0
transform 1 0 18906 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_353
timestamp 0
transform 1 0 19274 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_77_357
timestamp 0
transform 1 0 19458 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_359
timestamp 0
transform 1 0 19550 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_361
timestamp 0
transform 1 0 19642 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_369
timestamp 0
transform 1 0 20010 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_77_373
timestamp 0
transform 1 0 20194 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_77_381
timestamp 0
transform 1 0 20562 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_77_395
timestamp 0
transform 1 0 21206 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_403
timestamp 0
transform 1 0 21574 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_411
timestamp 0
transform 1 0 21942 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_77_419
timestamp 0
transform 1 0 22310 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_421
timestamp 0
transform 1 0 22402 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_77_429
timestamp 0
transform 1 0 22770 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_77_438
timestamp 0
transform 1 0 23184 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_77_447
timestamp 0
transform 1 0 23598 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_77_451
timestamp 0
transform 1 0 23782 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_453
timestamp 0
transform 1 0 23874 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_77_458
timestamp 0
transform 1 0 24104 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_77_465
timestamp 0
transform 1 0 24426 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_473
timestamp 0
transform 1 0 24794 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_77_477
timestamp 0
transform 1 0 24978 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_479
timestamp 0
transform 1 0 25070 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_481
timestamp 0
transform 1 0 25162 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_489
timestamp 0
transform 1 0 25530 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_497
timestamp 0
transform 1 0 25898 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_505
timestamp 0
transform 1 0 26266 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_513
timestamp 0
transform 1 0 26634 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_521
timestamp 0
transform 1 0 27002 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_529
timestamp 0
transform 1 0 27370 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_77_537
timestamp 0
transform 1 0 27738 0 -1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_77_539
timestamp 0
transform 1 0 27830 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_77_541
timestamp 0
transform 1 0 27922 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_549
timestamp 0
transform 1 0 28290 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_557
timestamp 0
transform 1 0 28658 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_565
timestamp 0
transform 1 0 29026 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_77_573
timestamp 0
transform 1 0 29394 0 -1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_77_581
timestamp 0
transform 1 0 29762 0 -1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_77_585
timestamp 0
transform 1 0 29946 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_78_0
timestamp 0
transform 1 0 3036 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_8
timestamp 0
transform 1 0 3404 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_16
timestamp 0
transform 1 0 3772 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_24
timestamp 0
transform 1 0 4140 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_28
timestamp 0
transform 1 0 4324 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_78_31
timestamp 0
transform 1 0 4462 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_39
timestamp 0
transform 1 0 4830 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_47
timestamp 0
transform 1 0 5198 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_51
timestamp 0
transform 1 0 5382 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_53
timestamp 0
transform 1 0 5474 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_78_78
timestamp 0
transform 1 0 6624 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_86
timestamp 0
transform 1 0 6992 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_91
timestamp 0
transform 1 0 7222 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_78_99
timestamp 0
transform 1 0 7590 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_101
timestamp 0
transform 1 0 7682 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_78_108
timestamp 0
transform 1 0 8004 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_136
timestamp 0
transform 1 0 9292 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_144
timestamp 0
transform 1 0 9660 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_148
timestamp 0
transform 1 0 9844 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_78_151
timestamp 0
transform 1 0 9982 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_78_159
timestamp 0
transform 1 0 10350 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_161
timestamp 0
transform 1 0 10442 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_78_170
timestamp 0
transform 1 0 10856 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_78_174
timestamp 0
transform 1 0 11040 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_78_199
timestamp 0
transform 1 0 12190 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_78_207
timestamp 0
transform 1 0 12558 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_209
timestamp 0
transform 1 0 12650 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_78_211
timestamp 0
transform 1 0 12742 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_215
timestamp 0
transform 1 0 12926 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_78_226
timestamp 0
transform 1 0 13432 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_243
timestamp 0
transform 1 0 14214 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_251
timestamp 0
transform 1 0 14582 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_78_264
timestamp 0
transform 1 0 15180 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_268
timestamp 0
transform 1 0 15364 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_78_271
timestamp 0
transform 1 0 15502 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_281
timestamp 0
transform 1 0 15962 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_289
timestamp 0
transform 1 0 16330 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_78_293
timestamp 0
transform 1 0 16514 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_78_311
timestamp 0
transform 1 0 17342 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_319
timestamp 0
transform 1 0 17710 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_78_327
timestamp 0
transform 1 0 18078 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_329
timestamp 0
transform 1 0 18170 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_78_331
timestamp 0
transform 1 0 18262 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_342
timestamp 0
transform 1 0 18768 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_350
timestamp 0
transform 1 0 19136 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_78_358
timestamp 0
transform 1 0 19504 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_78_383
timestamp 0
transform 1 0 20654 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_387
timestamp 0
transform 1 0 20838 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_389
timestamp 0
transform 1 0 20930 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_78_391
timestamp 0
transform 1 0 21022 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_399
timestamp 0
transform 1 0 21390 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_407
timestamp 0
transform 1 0 21758 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_435
timestamp 0
transform 1 0 23046 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_443
timestamp 0
transform 1 0 23414 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_447
timestamp 0
transform 1 0 23598 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_449
timestamp 0
transform 1 0 23690 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_78_451
timestamp 0
transform 1 0 23782 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_458
timestamp 0
transform 1 0 24104 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_466
timestamp 0
transform 1 0 24472 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_474
timestamp 0
transform 1 0 24840 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_482
timestamp 0
transform 1 0 25208 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_490
timestamp 0
transform 1 0 25576 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_498
timestamp 0
transform 1 0 25944 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_506
timestamp 0
transform 1 0 26312 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_78_511
timestamp 0
transform 1 0 26542 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_519
timestamp 0
transform 1 0 26910 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_527
timestamp 0
transform 1 0 27278 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_535
timestamp 0
transform 1 0 27646 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_543
timestamp 0
transform 1 0 28014 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_551
timestamp 0
transform 1 0 28382 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_78_559
timestamp 0
transform 1 0 28750 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_78_567
timestamp 0
transform 1 0 29118 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_569
timestamp 0
transform 1 0 29210 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_78_571
timestamp 0
transform 1 0 29302 0 1 24480
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_78_579
timestamp 0
transform 1 0 29670 0 1 24480
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_78_583
timestamp 0
transform 1 0 29854 0 1 24480
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_78_585
timestamp 0
transform 1 0 29946 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_79_0
timestamp 0
transform 1 0 3036 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_8
timestamp 0
transform 1 0 3404 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_16
timestamp 0
transform 1 0 3772 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_24
timestamp 0
transform 1 0 4140 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_32
timestamp 0
transform 1 0 4508 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_40
timestamp 0
transform 1 0 4876 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_48
timestamp 0
transform 1 0 5244 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_56
timestamp 0
transform 1 0 5612 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_79_61
timestamp 0
transform 1 0 5842 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_79_73
timestamp 0
transform 1 0 6394 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_81
timestamp 0
transform 1 0 6762 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_89
timestamp 0
transform 1 0 7130 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_97
timestamp 0
transform 1 0 7498 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_105
timestamp 0
transform 1 0 7866 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_113
timestamp 0
transform 1 0 8234 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_79_117
timestamp 0
transform 1 0 8418 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_79_119
timestamp 0
transform 1 0 8510 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_79_121
timestamp 0
transform 1 0 8602 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_129
timestamp 0
transform 1 0 8970 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_137
timestamp 0
transform 1 0 9338 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_79_141
timestamp 0
transform 1 0 9522 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_79_167
timestamp 0
transform 1 0 10718 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_175
timestamp 0
transform 1 0 11086 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_79_179
timestamp 0
transform 1 0 11270 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_79_181
timestamp 0
transform 1 0 11362 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_79_209
timestamp 0
transform 1 0 12650 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_79_226
timestamp 0
transform 1 0 13432 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_234
timestamp 0
transform 1 0 13800 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_79_238
timestamp 0
transform 1 0 13984 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_79_241
timestamp 0
transform 1 0 14122 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_249
timestamp 0
transform 1 0 14490 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_79_253
timestamp 0
transform 1 0 14674 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_79_255
timestamp 0
transform 1 0 14766 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_79_270
timestamp 0
transform 1 0 15456 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_79_274
timestamp 0
transform 1 0 15640 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_79_276
timestamp 0
transform 1 0 15732 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_79_283
timestamp 0
transform 1 0 16054 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_291
timestamp 0
transform 1 0 16422 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_79_299
timestamp 0
transform 1 0 16790 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_79_301
timestamp 0
transform 1 0 16882 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_79_314
timestamp 0
transform 1 0 17480 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_322
timestamp 0
transform 1 0 17848 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_79_330
timestamp 0
transform 1 0 18216 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_79_335
timestamp 0
transform 1 0 18446 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_79_346
timestamp 0
transform 1 0 18952 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_354
timestamp 0
transform 1 0 19320 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_79_358
timestamp 0
transform 1 0 19504 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_79_361
timestamp 0
transform 1 0 19642 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_369
timestamp 0
transform 1 0 20010 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_79_373
timestamp 0
transform 1 0 20194 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_79_381
timestamp 0
transform 1 0 20562 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_389
timestamp 0
transform 1 0 20930 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_404
timestamp 0
transform 1 0 21620 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_412
timestamp 0
transform 1 0 21988 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_421
timestamp 0
transform 1 0 22402 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_429
timestamp 0
transform 1 0 22770 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_437
timestamp 0
transform 1 0 23138 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_445
timestamp 0
transform 1 0 23506 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_453
timestamp 0
transform 1 0 23874 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_461
timestamp 0
transform 1 0 24242 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_469
timestamp 0
transform 1 0 24610 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_79_477
timestamp 0
transform 1 0 24978 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_79_479
timestamp 0
transform 1 0 25070 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_79_481
timestamp 0
transform 1 0 25162 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_489
timestamp 0
transform 1 0 25530 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_497
timestamp 0
transform 1 0 25898 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_505
timestamp 0
transform 1 0 26266 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_513
timestamp 0
transform 1 0 26634 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_521
timestamp 0
transform 1 0 27002 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_529
timestamp 0
transform 1 0 27370 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_79_537
timestamp 0
transform 1 0 27738 0 -1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_79_539
timestamp 0
transform 1 0 27830 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_79_541
timestamp 0
transform 1 0 27922 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_549
timestamp 0
transform 1 0 28290 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_557
timestamp 0
transform 1 0 28658 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_565
timestamp 0
transform 1 0 29026 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_79_573
timestamp 0
transform 1 0 29394 0 -1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_79_581
timestamp 0
transform 1 0 29762 0 -1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_79_585
timestamp 0
transform 1 0 29946 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_2  FILLER_80_0
timestamp 0
transform 1 0 3036 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_80_26
timestamp 0
transform 1 0 4232 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_80_31
timestamp 0
transform 1 0 4462 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_80_42
timestamp 0
transform 1 0 4968 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_50
timestamp 0
transform 1 0 5336 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_58
timestamp 0
transform 1 0 5704 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_66
timestamp 0
transform 1 0 6072 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_74
timestamp 0
transform 1 0 6440 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_82
timestamp 0
transform 1 0 6808 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_91
timestamp 0
transform 1 0 7222 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_99
timestamp 0
transform 1 0 7590 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_107
timestamp 0
transform 1 0 7958 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_115
timestamp 0
transform 1 0 8326 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_80_119
timestamp 0
transform 1 0 8510 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_80_121
timestamp 0
transform 1 0 8602 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_80_146
timestamp 0
transform 1 0 9752 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_80_151
timestamp 0
transform 1 0 9982 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_159
timestamp 0
transform 1 0 10350 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_167
timestamp 0
transform 1 0 10718 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_80_171
timestamp 0
transform 1 0 10902 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_80_197
timestamp 0
transform 1 0 12098 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_205
timestamp 0
transform 1 0 12466 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_80_209
timestamp 0
transform 1 0 12650 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_80_211
timestamp 0
transform 1 0 12742 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_219
timestamp 0
transform 1 0 13110 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_227
timestamp 0
transform 1 0 13478 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_235
timestamp 0
transform 1 0 13846 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_243
timestamp 0
transform 1 0 14214 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_251
timestamp 0
transform 1 0 14582 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_80_255
timestamp 0
transform 1 0 14766 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_80_262
timestamp 0
transform 1 0 15088 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_271
timestamp 0
transform 1 0 15502 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_279
timestamp 0
transform 1 0 15870 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_287
timestamp 0
transform 1 0 16238 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_295
timestamp 0
transform 1 0 16606 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_80_303
timestamp 0
transform 1 0 16974 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_80_305
timestamp 0
transform 1 0 17066 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_80_313
timestamp 0
transform 1 0 17434 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_80_321
timestamp 0
transform 1 0 17802 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_80_329
timestamp 0
transform 1 0 18170 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_80_331
timestamp 0
transform 1 0 18262 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_80_335
timestamp 0
transform 1 0 18446 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_80_352
timestamp 0
transform 1 0 19228 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_360
timestamp 0
transform 1 0 19596 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_368
timestamp 0
transform 1 0 19964 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_80_372
timestamp 0
transform 1 0 20148 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_80_381
timestamp 0
transform 1 0 20562 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_80_389
timestamp 0
transform 1 0 20930 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_80_391
timestamp 0
transform 1 0 21022 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_399
timestamp 0
transform 1 0 21390 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_80_403
timestamp 0
transform 1 0 21574 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_80_429
timestamp 0
transform 1 0 22770 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_437
timestamp 0
transform 1 0 23138 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_445
timestamp 0
transform 1 0 23506 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_80_449
timestamp 0
transform 1 0 23690 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_80_451
timestamp 0
transform 1 0 23782 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_459
timestamp 0
transform 1 0 24150 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_467
timestamp 0
transform 1 0 24518 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_475
timestamp 0
transform 1 0 24886 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_483
timestamp 0
transform 1 0 25254 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_491
timestamp 0
transform 1 0 25622 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_499
timestamp 0
transform 1 0 25990 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_80_507
timestamp 0
transform 1 0 26358 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_80_509
timestamp 0
transform 1 0 26450 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_80_511
timestamp 0
transform 1 0 26542 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_519
timestamp 0
transform 1 0 26910 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_527
timestamp 0
transform 1 0 27278 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_535
timestamp 0
transform 1 0 27646 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_543
timestamp 0
transform 1 0 28014 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_551
timestamp 0
transform 1 0 28382 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_80_559
timestamp 0
transform 1 0 28750 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_80_567
timestamp 0
transform 1 0 29118 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_80_569
timestamp 0
transform 1 0 29210 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_80_571
timestamp 0
transform 1 0 29302 0 1 25024
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_80_579
timestamp 0
transform 1 0 29670 0 1 25024
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_80_583
timestamp 0
transform 1 0 29854 0 1 25024
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_80_585
timestamp 0
transform 1 0 29946 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_81_0
timestamp 0
transform 1 0 3036 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_81_4
timestamp 0
transform 1 0 3220 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_6
timestamp 0
transform 1 0 3312 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_31
timestamp 0
transform 1 0 4462 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_39
timestamp 0
transform 1 0 4830 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_47
timestamp 0
transform 1 0 5198 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_55
timestamp 0
transform 1 0 5566 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_81_59
timestamp 0
transform 1 0 5750 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_61
timestamp 0
transform 1 0 5842 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_69
timestamp 0
transform 1 0 6210 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_81_73
timestamp 0
transform 1 0 6394 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_81_99
timestamp 0
transform 1 0 7590 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_81_107
timestamp 0
transform 1 0 7958 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_81_113
timestamp 0
transform 1 0 8234 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_81_117
timestamp 0
transform 1 0 8418 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_119
timestamp 0
transform 1 0 8510 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_121
timestamp 0
transform 1 0 8602 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_129
timestamp 0
transform 1 0 8970 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_137
timestamp 0
transform 1 0 9338 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_81_141
timestamp 0
transform 1 0 9522 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_143
timestamp 0
transform 1 0 9614 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_168
timestamp 0
transform 1 0 10764 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_176
timestamp 0
transform 1 0 11132 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_81_181
timestamp 0
transform 1 0 11362 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_189
timestamp 0
transform 1 0 11730 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_197
timestamp 0
transform 1 0 12098 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_205
timestamp 0
transform 1 0 12466 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_213
timestamp 0
transform 1 0 12834 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_221
timestamp 0
transform 1 0 13202 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_229
timestamp 0
transform 1 0 13570 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_81_237
timestamp 0
transform 1 0 13938 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_239
timestamp 0
transform 1 0 14030 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_241
timestamp 0
transform 1 0 14122 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_249
timestamp 0
transform 1 0 14490 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_257
timestamp 0
transform 1 0 14858 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_265
timestamp 0
transform 1 0 15226 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_273
timestamp 0
transform 1 0 15594 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_281
timestamp 0
transform 1 0 15962 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_289
timestamp 0
transform 1 0 16330 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_81_297
timestamp 0
transform 1 0 16698 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_299
timestamp 0
transform 1 0 16790 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_301
timestamp 0
transform 1 0 16882 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_309
timestamp 0
transform 1 0 17250 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_317
timestamp 0
transform 1 0 17618 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_325
timestamp 0
transform 1 0 17986 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_333
timestamp 0
transform 1 0 18354 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_81_337
timestamp 0
transform 1 0 18538 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_81_345
timestamp 0
transform 1 0 18906 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_81_353
timestamp 0
transform 1 0 19274 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_81_357
timestamp 0
transform 1 0 19458 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_359
timestamp 0
transform 1 0 19550 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_361
timestamp 0
transform 1 0 19642 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_369
timestamp 0
transform 1 0 20010 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_377
timestamp 0
transform 1 0 20378 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_385
timestamp 0
transform 1 0 20746 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_393
timestamp 0
transform 1 0 21114 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_401
timestamp 0
transform 1 0 21482 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_409
timestamp 0
transform 1 0 21850 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_81_417
timestamp 0
transform 1 0 22218 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_419
timestamp 0
transform 1 0 22310 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_421
timestamp 0
transform 1 0 22402 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_429
timestamp 0
transform 1 0 22770 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_437
timestamp 0
transform 1 0 23138 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_81_441
timestamp 0
transform 1 0 23322 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_81_450
timestamp 0
transform 1 0 23736 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_458
timestamp 0
transform 1 0 24104 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_466
timestamp 0
transform 1 0 24472 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_474
timestamp 0
transform 1 0 24840 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_81_478
timestamp 0
transform 1 0 25024 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_81_481
timestamp 0
transform 1 0 25162 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_489
timestamp 0
transform 1 0 25530 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_497
timestamp 0
transform 1 0 25898 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_505
timestamp 0
transform 1 0 26266 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_513
timestamp 0
transform 1 0 26634 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_521
timestamp 0
transform 1 0 27002 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_529
timestamp 0
transform 1 0 27370 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_81_537
timestamp 0
transform 1 0 27738 0 -1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_81_539
timestamp 0
transform 1 0 27830 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_81_541
timestamp 0
transform 1 0 27922 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_549
timestamp 0
transform 1 0 28290 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_557
timestamp 0
transform 1 0 28658 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_565
timestamp 0
transform 1 0 29026 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_81_573
timestamp 0
transform 1 0 29394 0 -1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_81_581
timestamp 0
transform 1 0 29762 0 -1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_81_585
timestamp 0
transform 1 0 29946 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_0
timestamp 0
transform 1 0 3036 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_8
timestamp 0
transform 1 0 3404 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_16
timestamp 0
transform 1 0 3772 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_24
timestamp 0
transform 1 0 4140 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_82_28
timestamp 0
transform 1 0 4324 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_82_31
timestamp 0
transform 1 0 4462 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_82_59
timestamp 0
transform 1 0 5750 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_67
timestamp 0
transform 1 0 6118 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_75
timestamp 0
transform 1 0 6486 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_83
timestamp 0
transform 1 0 6854 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_82_87
timestamp 0
transform 1 0 7038 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_82_89
timestamp 0
transform 1 0 7130 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_91
timestamp 0
transform 1 0 7222 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_82_99
timestamp 0
transform 1 0 7590 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_82_101
timestamp 0
transform 1 0 7682 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_82_105
timestamp 0
transform 1 0 7866 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_82_109
timestamp 0
transform 1 0 8050 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_82_125
timestamp 0
transform 1 0 8786 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_82_134
timestamp 0
transform 1 0 9200 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_142
timestamp 0
transform 1 0 9568 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_151
timestamp 0
transform 1 0 9982 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_159
timestamp 0
transform 1 0 10350 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_167
timestamp 0
transform 1 0 10718 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_175
timestamp 0
transform 1 0 11086 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_183
timestamp 0
transform 1 0 11454 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_191
timestamp 0
transform 1 0 11822 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_199
timestamp 0
transform 1 0 12190 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_82_207
timestamp 0
transform 1 0 12558 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_82_209
timestamp 0
transform 1 0 12650 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_211
timestamp 0
transform 1 0 12742 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_219
timestamp 0
transform 1 0 13110 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_227
timestamp 0
transform 1 0 13478 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_82_234
timestamp 0
transform 1 0 13800 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_242
timestamp 0
transform 1 0 14168 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_250
timestamp 0
transform 1 0 14536 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_258
timestamp 0
transform 1 0 14904 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_266
timestamp 0
transform 1 0 15272 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_82_271
timestamp 0
transform 1 0 15502 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_279
timestamp 0
transform 1 0 15870 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_82_283
timestamp 0
transform 1 0 16054 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_291
timestamp 0
transform 1 0 16422 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_299
timestamp 0
transform 1 0 16790 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 0
transform 1 0 17158 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_315
timestamp 0
transform 1 0 17526 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_323
timestamp 0
transform 1 0 17894 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_82_327
timestamp 0
transform 1 0 18078 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_82_329
timestamp 0
transform 1 0 18170 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_331
timestamp 0
transform 1 0 18262 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_339
timestamp 0
transform 1 0 18630 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_347
timestamp 0
transform 1 0 18998 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_355
timestamp 0
transform 1 0 19366 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_363
timestamp 0
transform 1 0 19734 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_371
timestamp 0
transform 1 0 20102 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_82_379
timestamp 0
transform 1 0 20470 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_82_384
timestamp 0
transform 1 0 20700 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_82_388
timestamp 0
transform 1 0 20884 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_82_391
timestamp 0
transform 1 0 21022 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_399
timestamp 0
transform 1 0 21390 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_82_406
timestamp 0
transform 1 0 21712 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_414
timestamp 0
transform 1 0 22080 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_422
timestamp 0
transform 1 0 22448 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_437
timestamp 0
transform 1 0 23138 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_445
timestamp 0
transform 1 0 23506 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_82_449
timestamp 0
transform 1 0 23690 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_451
timestamp 0
transform 1 0 23782 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_459
timestamp 0
transform 1 0 24150 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_467
timestamp 0
transform 1 0 24518 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_475
timestamp 0
transform 1 0 24886 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_483
timestamp 0
transform 1 0 25254 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_491
timestamp 0
transform 1 0 25622 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_499
timestamp 0
transform 1 0 25990 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_82_507
timestamp 0
transform 1 0 26358 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_82_509
timestamp 0
transform 1 0 26450 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_511
timestamp 0
transform 1 0 26542 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_519
timestamp 0
transform 1 0 26910 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_527
timestamp 0
transform 1 0 27278 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_535
timestamp 0
transform 1 0 27646 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_543
timestamp 0
transform 1 0 28014 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_551
timestamp 0
transform 1 0 28382 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_82_559
timestamp 0
transform 1 0 28750 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_82_567
timestamp 0
transform 1 0 29118 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_82_569
timestamp 0
transform 1 0 29210 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_82_571
timestamp 0
transform 1 0 29302 0 1 25568
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_82_579
timestamp 0
transform 1 0 29670 0 1 25568
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_82_583
timestamp 0
transform 1 0 29854 0 1 25568
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_82_585
timestamp 0
transform 1 0 29946 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_83_0
timestamp 0
transform 1 0 3036 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_8
timestamp 0
transform 1 0 3404 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_16
timestamp 0
transform 1 0 3772 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_24
timestamp 0
transform 1 0 4140 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_83_28
timestamp 0
transform 1 0 4324 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_83_54
timestamp 0
transform 1 0 5520 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_83_58
timestamp 0
transform 1 0 5704 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_83_61
timestamp 0
transform 1 0 5842 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_69
timestamp 0
transform 1 0 6210 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_83_77
timestamp 0
transform 1 0 6578 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_83_88
timestamp 0
transform 1 0 7084 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_83_116
timestamp 0
transform 1 0 8372 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_83_121
timestamp 0
transform 1 0 8602 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_83_129
timestamp 0
transform 1 0 8970 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_83_155
timestamp 0
transform 1 0 10166 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_163
timestamp 0
transform 1 0 10534 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_171
timestamp 0
transform 1 0 10902 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_83_179
timestamp 0
transform 1 0 11270 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_83_181
timestamp 0
transform 1 0 11362 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_189
timestamp 0
transform 1 0 11730 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_197
timestamp 0
transform 1 0 12098 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_205
timestamp 0
transform 1 0 12466 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_83_213
timestamp 0
transform 1 0 12834 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_83_226
timestamp 0
transform 1 0 13432 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_83_234
timestamp 0
transform 1 0 13800 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_83_238
timestamp 0
transform 1 0 13984 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_83_241
timestamp 0
transform 1 0 14122 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_249
timestamp 0
transform 1 0 14490 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_257
timestamp 0
transform 1 0 14858 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_265
timestamp 0
transform 1 0 15226 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_273
timestamp 0
transform 1 0 15594 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_281
timestamp 0
transform 1 0 15962 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_289
timestamp 0
transform 1 0 16330 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_83_297
timestamp 0
transform 1 0 16698 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_83_299
timestamp 0
transform 1 0 16790 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_83_301
timestamp 0
transform 1 0 16882 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_309
timestamp 0
transform 1 0 17250 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_317
timestamp 0
transform 1 0 17618 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_83_337
timestamp 0
transform 1 0 18538 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_345
timestamp 0
transform 1 0 18906 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_353
timestamp 0
transform 1 0 19274 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_83_357
timestamp 0
transform 1 0 19458 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_83_359
timestamp 0
transform 1 0 19550 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_83_361
timestamp 0
transform 1 0 19642 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_369
timestamp 0
transform 1 0 20010 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_83_397
timestamp 0
transform 1 0 21298 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_83_406
timestamp 0
transform 1 0 21712 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_414
timestamp 0
transform 1 0 22080 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_83_418
timestamp 0
transform 1 0 22264 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_83_421
timestamp 0
transform 1 0 22402 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_429
timestamp 0
transform 1 0 22770 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_83_433
timestamp 0
transform 1 0 22954 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_83_435
timestamp 0
transform 1 0 23046 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_83_443
timestamp 0
transform 1 0 23414 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_451
timestamp 0
transform 1 0 23782 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_459
timestamp 0
transform 1 0 24150 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_467
timestamp 0
transform 1 0 24518 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_475
timestamp 0
transform 1 0 24886 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_83_479
timestamp 0
transform 1 0 25070 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_83_481
timestamp 0
transform 1 0 25162 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_489
timestamp 0
transform 1 0 25530 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_497
timestamp 0
transform 1 0 25898 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_505
timestamp 0
transform 1 0 26266 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_513
timestamp 0
transform 1 0 26634 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_521
timestamp 0
transform 1 0 27002 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_529
timestamp 0
transform 1 0 27370 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_83_537
timestamp 0
transform 1 0 27738 0 -1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_83_539
timestamp 0
transform 1 0 27830 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_83_541
timestamp 0
transform 1 0 27922 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_549
timestamp 0
transform 1 0 28290 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_557
timestamp 0
transform 1 0 28658 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_565
timestamp 0
transform 1 0 29026 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_83_573
timestamp 0
transform 1 0 29394 0 -1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_83_581
timestamp 0
transform 1 0 29762 0 -1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_83_585
timestamp 0
transform 1 0 29946 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_0
timestamp 0
transform 1 0 3036 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_8
timestamp 0
transform 1 0 3404 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_16
timestamp 0
transform 1 0 3772 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_84_24
timestamp 0
transform 1 0 4140 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_84_28
timestamp 0
transform 1 0 4324 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_84_31
timestamp 0
transform 1 0 4462 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_39
timestamp 0
transform 1 0 4830 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_84_47
timestamp 0
transform 1 0 5198 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_84_51
timestamp 0
transform 1 0 5382 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_53
timestamp 0
transform 1 0 5474 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_78
timestamp 0
transform 1 0 6624 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_84_86
timestamp 0
transform 1 0 6992 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_84_91
timestamp 0
transform 1 0 7222 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_84_99
timestamp 0
transform 1 0 7590 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_84_112
timestamp 0
transform 1 0 8188 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_84_116
timestamp 0
transform 1 0 8372 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_141
timestamp 0
transform 1 0 9522 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_84_149
timestamp 0
transform 1 0 9890 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_151
timestamp 0
transform 1 0 9982 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_159
timestamp 0
transform 1 0 10350 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_167
timestamp 0
transform 1 0 10718 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_175
timestamp 0
transform 1 0 11086 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_84_183
timestamp 0
transform 1 0 11454 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_185
timestamp 0
transform 1 0 11546 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_189
timestamp 0
transform 1 0 11730 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_200
timestamp 0
transform 1 0 12236 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_84_208
timestamp 0
transform 1 0 12604 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_84_211
timestamp 0
transform 1 0 12742 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_84_226
timestamp 0
transform 1 0 13432 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_84_246
timestamp 0
transform 1 0 14352 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_84_254
timestamp 0
transform 1 0 14720 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_84_264
timestamp 0
transform 1 0 15180 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_84_268
timestamp 0
transform 1 0 15364 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_84_271
timestamp 0
transform 1 0 15502 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_84_279
timestamp 0
transform 1 0 15870 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_84_283
timestamp 0
transform 1 0 16054 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_285
timestamp 0
transform 1 0 16146 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_292
timestamp 0
transform 1 0 16468 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_300
timestamp 0
transform 1 0 16836 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_308
timestamp 0
transform 1 0 17204 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_84_316
timestamp 0
transform 1 0 17572 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_318
timestamp 0
transform 1 0 17664 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_84_325
timestamp 0
transform 1 0 17986 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_84_329
timestamp 0
transform 1 0 18170 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_331
timestamp 0
transform 1 0 18262 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_339
timestamp 0
transform 1 0 18630 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_84_347
timestamp 0
transform 1 0 18998 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_84_373
timestamp 0
transform 1 0 20194 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_381
timestamp 0
transform 1 0 20562 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_84_389
timestamp 0
transform 1 0 20930 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_391
timestamp 0
transform 1 0 21022 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_399
timestamp 0
transform 1 0 21390 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_407
timestamp 0
transform 1 0 21758 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_415
timestamp 0
transform 1 0 22126 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_423
timestamp 0
transform 1 0 22494 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_431
timestamp 0
transform 1 0 22862 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_439
timestamp 0
transform 1 0 23230 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_84_447
timestamp 0
transform 1 0 23598 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_449
timestamp 0
transform 1 0 23690 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_451
timestamp 0
transform 1 0 23782 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_459
timestamp 0
transform 1 0 24150 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_467
timestamp 0
transform 1 0 24518 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_475
timestamp 0
transform 1 0 24886 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_483
timestamp 0
transform 1 0 25254 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_491
timestamp 0
transform 1 0 25622 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_499
timestamp 0
transform 1 0 25990 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_84_507
timestamp 0
transform 1 0 26358 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_509
timestamp 0
transform 1 0 26450 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_511
timestamp 0
transform 1 0 26542 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_519
timestamp 0
transform 1 0 26910 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_527
timestamp 0
transform 1 0 27278 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_535
timestamp 0
transform 1 0 27646 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_543
timestamp 0
transform 1 0 28014 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_551
timestamp 0
transform 1 0 28382 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_84_559
timestamp 0
transform 1 0 28750 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_84_567
timestamp 0
transform 1 0 29118 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_569
timestamp 0
transform 1 0 29210 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_84_571
timestamp 0
transform 1 0 29302 0 1 26112
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_84_579
timestamp 0
transform 1 0 29670 0 1 26112
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_84_583
timestamp 0
transform 1 0 29854 0 1 26112
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_84_585
timestamp 0
transform 1 0 29946 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_85_0
timestamp 0
transform 1 0 3036 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_8
timestamp 0
transform 1 0 3404 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_16
timestamp 0
transform 1 0 3772 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_24
timestamp 0
transform 1 0 4140 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_32
timestamp 0
transform 1 0 4508 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_40
timestamp 0
transform 1 0 4876 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_48
timestamp 0
transform 1 0 5244 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_56
timestamp 0
transform 1 0 5612 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_85_61
timestamp 0
transform 1 0 5842 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_85_74
timestamp 0
transform 1 0 6440 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_85_82
timestamp 0
transform 1 0 6808 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_85_94
timestamp 0
transform 1 0 7360 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_102
timestamp 0
transform 1 0 7728 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_110
timestamp 0
transform 1 0 8096 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_85_118
timestamp 0
transform 1 0 8464 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_85_121
timestamp 0
transform 1 0 8602 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_85_129
timestamp 0
transform 1 0 8970 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_85_140
timestamp 0
transform 1 0 9476 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_148
timestamp 0
transform 1 0 9844 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_156
timestamp 0
transform 1 0 10212 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_85_160
timestamp 0
transform 1 0 10396 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_85_168
timestamp 0
transform 1 0 10764 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_176
timestamp 0
transform 1 0 11132 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_85_181
timestamp 0
transform 1 0 11362 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_205
timestamp 0
transform 1 0 12466 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_213
timestamp 0
transform 1 0 12834 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_221
timestamp 0
transform 1 0 13202 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_85_225
timestamp 0
transform 1 0 13386 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_85_232
timestamp 0
transform 1 0 13708 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_241
timestamp 0
transform 1 0 14122 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_249
timestamp 0
transform 1 0 14490 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_257
timestamp 0
transform 1 0 14858 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_85_261
timestamp 0
transform 1 0 15042 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_85_269
timestamp 0
transform 1 0 15410 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_281
timestamp 0
transform 1 0 15962 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_85_292
timestamp 0
transform 1 0 16468 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_301
timestamp 0
transform 1 0 16882 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_309
timestamp 0
transform 1 0 17250 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_85_317
timestamp 0
transform 1 0 17618 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_85_326
timestamp 0
transform 1 0 18032 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_85_333
timestamp 0
transform 1 0 18354 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_341
timestamp 0
transform 1 0 18722 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_349
timestamp 0
transform 1 0 19090 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_85_357
timestamp 0
transform 1 0 19458 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_85_359
timestamp 0
transform 1 0 19550 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_85_361
timestamp 0
transform 1 0 19642 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_369
timestamp 0
transform 1 0 20010 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_386
timestamp 0
transform 1 0 20792 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_85_390
timestamp 0
transform 1 0 20976 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_85_416
timestamp 0
transform 1 0 22172 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_85_421
timestamp 0
transform 1 0 22402 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_429
timestamp 0
transform 1 0 22770 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_437
timestamp 0
transform 1 0 23138 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_445
timestamp 0
transform 1 0 23506 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_453
timestamp 0
transform 1 0 23874 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_461
timestamp 0
transform 1 0 24242 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_469
timestamp 0
transform 1 0 24610 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_85_477
timestamp 0
transform 1 0 24978 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_85_479
timestamp 0
transform 1 0 25070 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_85_481
timestamp 0
transform 1 0 25162 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_489
timestamp 0
transform 1 0 25530 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_497
timestamp 0
transform 1 0 25898 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_505
timestamp 0
transform 1 0 26266 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_513
timestamp 0
transform 1 0 26634 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_521
timestamp 0
transform 1 0 27002 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_529
timestamp 0
transform 1 0 27370 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_85_537
timestamp 0
transform 1 0 27738 0 -1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_85_539
timestamp 0
transform 1 0 27830 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_85_541
timestamp 0
transform 1 0 27922 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_549
timestamp 0
transform 1 0 28290 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_557
timestamp 0
transform 1 0 28658 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_565
timestamp 0
transform 1 0 29026 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_85_573
timestamp 0
transform 1 0 29394 0 -1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_85_581
timestamp 0
transform 1 0 29762 0 -1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_85_585
timestamp 0
transform 1 0 29946 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_86_0
timestamp 0
transform 1 0 3036 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_8
timestamp 0
transform 1 0 3404 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_16
timestamp 0
transform 1 0 3772 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_86_24
timestamp 0
transform 1 0 4140 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_86_28
timestamp 0
transform 1 0 4324 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_86_31
timestamp 0
transform 1 0 4462 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_39
timestamp 0
transform 1 0 4830 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_47
timestamp 0
transform 1 0 5198 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_55
timestamp 0
transform 1 0 5566 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_63
timestamp 0
transform 1 0 5934 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_86_71
timestamp 0
transform 1 0 6302 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_86_86
timestamp 0
transform 1 0 6992 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_86_91
timestamp 0
transform 1 0 7222 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_86_102
timestamp 0
transform 1 0 7728 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_86_110
timestamp 0
transform 1 0 8096 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_86_114
timestamp 0
transform 1 0 8280 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_86_124
timestamp 0
transform 1 0 8740 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_132
timestamp 0
transform 1 0 9108 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_140
timestamp 0
transform 1 0 9476 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_86_148
timestamp 0
transform 1 0 9844 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_86_151
timestamp 0
transform 1 0 9982 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_86_155
timestamp 0
transform 1 0 10166 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_86_173
timestamp 0
transform 1 0 10994 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_86_177
timestamp 0
transform 1 0 11178 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_86_195
timestamp 0
transform 1 0 12006 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_86_202
timestamp 0
transform 1 0 12328 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_211
timestamp 0
transform 1 0 12742 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_219
timestamp 0
transform 1 0 13110 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_227
timestamp 0
transform 1 0 13478 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_235
timestamp 0
transform 1 0 13846 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_243
timestamp 0
transform 1 0 14214 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_86_253
timestamp 0
transform 1 0 14674 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_86_262
timestamp 0
transform 1 0 15088 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_271
timestamp 0
transform 1 0 15502 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_279
timestamp 0
transform 1 0 15870 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_86_287
timestamp 0
transform 1 0 16238 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_86_291
timestamp 0
transform 1 0 16422 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_86_308
timestamp 0
transform 1 0 17204 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_86_316
timestamp 0
transform 1 0 17572 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_86_320
timestamp 0
transform 1 0 17756 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_86_326
timestamp 0
transform 1 0 18032 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_86_331
timestamp 0
transform 1 0 18262 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_339
timestamp 0
transform 1 0 18630 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_86_347
timestamp 0
transform 1 0 18998 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_86_349
timestamp 0
transform 1 0 19090 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_86_374
timestamp 0
transform 1 0 20240 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_382
timestamp 0
transform 1 0 20608 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_391
timestamp 0
transform 1 0 21022 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_399
timestamp 0
transform 1 0 21390 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_407
timestamp 0
transform 1 0 21758 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_415
timestamp 0
transform 1 0 22126 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_423
timestamp 0
transform 1 0 22494 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_431
timestamp 0
transform 1 0 22862 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_439
timestamp 0
transform 1 0 23230 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_86_447
timestamp 0
transform 1 0 23598 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_86_449
timestamp 0
transform 1 0 23690 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_86_451
timestamp 0
transform 1 0 23782 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_459
timestamp 0
transform 1 0 24150 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_467
timestamp 0
transform 1 0 24518 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_475
timestamp 0
transform 1 0 24886 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_483
timestamp 0
transform 1 0 25254 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_491
timestamp 0
transform 1 0 25622 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_499
timestamp 0
transform 1 0 25990 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_86_507
timestamp 0
transform 1 0 26358 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_86_509
timestamp 0
transform 1 0 26450 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_86_511
timestamp 0
transform 1 0 26542 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_519
timestamp 0
transform 1 0 26910 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_527
timestamp 0
transform 1 0 27278 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_535
timestamp 0
transform 1 0 27646 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_543
timestamp 0
transform 1 0 28014 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_551
timestamp 0
transform 1 0 28382 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_86_559
timestamp 0
transform 1 0 28750 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_86_567
timestamp 0
transform 1 0 29118 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_86_569
timestamp 0
transform 1 0 29210 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_86_571
timestamp 0
transform 1 0 29302 0 1 26656
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_86_579
timestamp 0
transform 1 0 29670 0 1 26656
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_86_583
timestamp 0
transform 1 0 29854 0 1 26656
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_86_585
timestamp 0
transform 1 0 29946 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_87_0
timestamp 0
transform 1 0 3036 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_8
timestamp 0
transform 1 0 3404 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_16
timestamp 0
transform 1 0 3772 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_24
timestamp 0
transform 1 0 4140 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_56
timestamp 0
transform 1 0 5612 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_87_61
timestamp 0
transform 1 0 5842 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_87_74
timestamp 0
transform 1 0 6440 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_87_78
timestamp 0
transform 1 0 6624 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_87_104
timestamp 0
transform 1 0 7820 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_87_108
timestamp 0
transform 1 0 8004 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_87_110
timestamp 0
transform 1 0 8096 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_87_116
timestamp 0
transform 1 0 8372 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_87_121
timestamp 0
transform 1 0 8602 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_87_131
timestamp 0
transform 1 0 9062 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_87_139
timestamp 0
transform 1 0 9430 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_147
timestamp 0
transform 1 0 9798 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_155
timestamp 0
transform 1 0 10166 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_87_163
timestamp 0
transform 1 0 10534 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_87_170
timestamp 0
transform 1 0 10856 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_87_178
timestamp 0
transform 1 0 11224 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_87_181
timestamp 0
transform 1 0 11362 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_87_189
timestamp 0
transform 1 0 11730 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_87_195
timestamp 0
transform 1 0 12006 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_87_202
timestamp 0
transform 1 0 12328 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_210
timestamp 0
transform 1 0 12696 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_218
timestamp 0
transform 1 0 13064 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_87_222
timestamp 0
transform 1 0 13248 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_87_228
timestamp 0
transform 1 0 13524 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_236
timestamp 0
transform 1 0 13892 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_87_241
timestamp 0
transform 1 0 14122 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_87_249
timestamp 0
transform 1 0 14490 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_87_267
timestamp 0
transform 1 0 15318 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_275
timestamp 0
transform 1 0 15686 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_283
timestamp 0
transform 1 0 16054 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_87_287
timestamp 0
transform 1 0 16238 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_87_295
timestamp 0
transform 1 0 16606 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_87_299
timestamp 0
transform 1 0 16790 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_87_301
timestamp 0
transform 1 0 16882 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_309
timestamp 0
transform 1 0 17250 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_317
timestamp 0
transform 1 0 17618 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_325
timestamp 0
transform 1 0 17986 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_87_329
timestamp 0
transform 1 0 18170 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_87_334
timestamp 0
transform 1 0 18400 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_342
timestamp 0
transform 1 0 18768 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_350
timestamp 0
transform 1 0 19136 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_87_358
timestamp 0
transform 1 0 19504 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_87_361
timestamp 0
transform 1 0 19642 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_369
timestamp 0
transform 1 0 20010 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_87_373
timestamp 0
transform 1 0 20194 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_87_398
timestamp 0
transform 1 0 21344 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_406
timestamp 0
transform 1 0 21712 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_414
timestamp 0
transform 1 0 22080 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_87_418
timestamp 0
transform 1 0 22264 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_87_421
timestamp 0
transform 1 0 22402 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_429
timestamp 0
transform 1 0 22770 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_437
timestamp 0
transform 1 0 23138 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_445
timestamp 0
transform 1 0 23506 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_453
timestamp 0
transform 1 0 23874 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_461
timestamp 0
transform 1 0 24242 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_469
timestamp 0
transform 1 0 24610 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_87_477
timestamp 0
transform 1 0 24978 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_87_479
timestamp 0
transform 1 0 25070 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_87_481
timestamp 0
transform 1 0 25162 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_489
timestamp 0
transform 1 0 25530 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_497
timestamp 0
transform 1 0 25898 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_505
timestamp 0
transform 1 0 26266 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_513
timestamp 0
transform 1 0 26634 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_521
timestamp 0
transform 1 0 27002 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_529
timestamp 0
transform 1 0 27370 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_87_537
timestamp 0
transform 1 0 27738 0 -1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_87_539
timestamp 0
transform 1 0 27830 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_87_541
timestamp 0
transform 1 0 27922 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_549
timestamp 0
transform 1 0 28290 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_557
timestamp 0
transform 1 0 28658 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_565
timestamp 0
transform 1 0 29026 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_87_573
timestamp 0
transform 1 0 29394 0 -1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_87_581
timestamp 0
transform 1 0 29762 0 -1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_87_585
timestamp 0
transform 1 0 29946 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_0
timestamp 0
transform 1 0 3036 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_8
timestamp 0
transform 1 0 3404 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_16
timestamp 0
transform 1 0 3772 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_88_24
timestamp 0
transform 1 0 4140 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_88_28
timestamp 0
transform 1 0 4324 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_88_31
timestamp 0
transform 1 0 4462 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_39
timestamp 0
transform 1 0 4830 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_88_47
timestamp 0
transform 1 0 5198 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_49
timestamp 0
transform 1 0 5290 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_74
timestamp 0
transform 1 0 6440 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_82
timestamp 0
transform 1 0 6808 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_88_91
timestamp 0
transform 1 0 7222 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_88_102
timestamp 0
transform 1 0 7728 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_110
timestamp 0
transform 1 0 8096 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_88_118
timestamp 0
transform 1 0 8464 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_120
timestamp 0
transform 1 0 8556 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_88_128
timestamp 0
transform 1 0 8924 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_88_132
timestamp 0
transform 1 0 9108 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_134
timestamp 0
transform 1 0 9200 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_88_146
timestamp 0
transform 1 0 9752 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_88_151
timestamp 0
transform 1 0 9982 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_159
timestamp 0
transform 1 0 10350 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_167
timestamp 0
transform 1 0 10718 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_175
timestamp 0
transform 1 0 11086 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_183
timestamp 0
transform 1 0 11454 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_191
timestamp 0
transform 1 0 11822 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_199
timestamp 0
transform 1 0 12190 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_88_207
timestamp 0
transform 1 0 12558 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_209
timestamp 0
transform 1 0 12650 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_211
timestamp 0
transform 1 0 12742 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_235
timestamp 0
transform 1 0 13846 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_243
timestamp 0
transform 1 0 14214 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_251
timestamp 0
transform 1 0 14582 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_88_263
timestamp 0
transform 1 0 15134 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_88_267
timestamp 0
transform 1 0 15318 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_269
timestamp 0
transform 1 0 15410 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_271
timestamp 0
transform 1 0 15502 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_279
timestamp 0
transform 1 0 15870 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_88_287
timestamp 0
transform 1 0 16238 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_88_291
timestamp 0
transform 1 0 16422 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_295
timestamp 0
transform 1 0 16606 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_303
timestamp 0
transform 1 0 16974 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_311
timestamp 0
transform 1 0 17342 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_319
timestamp 0
transform 1 0 17710 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_88_327
timestamp 0
transform 1 0 18078 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_329
timestamp 0
transform 1 0 18170 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_331
timestamp 0
transform 1 0 18262 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_88_343
timestamp 0
transform 1 0 18814 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_88_347
timestamp 0
transform 1 0 18998 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_349
timestamp 0
transform 1 0 19090 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_374
timestamp 0
transform 1 0 20240 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_382
timestamp 0
transform 1 0 20608 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_391
timestamp 0
transform 1 0 21022 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_399
timestamp 0
transform 1 0 21390 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_407
timestamp 0
transform 1 0 21758 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_415
timestamp 0
transform 1 0 22126 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_423
timestamp 0
transform 1 0 22494 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_431
timestamp 0
transform 1 0 22862 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_439
timestamp 0
transform 1 0 23230 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_88_447
timestamp 0
transform 1 0 23598 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_449
timestamp 0
transform 1 0 23690 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_451
timestamp 0
transform 1 0 23782 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_459
timestamp 0
transform 1 0 24150 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_467
timestamp 0
transform 1 0 24518 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_475
timestamp 0
transform 1 0 24886 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_483
timestamp 0
transform 1 0 25254 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_491
timestamp 0
transform 1 0 25622 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_499
timestamp 0
transform 1 0 25990 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_88_507
timestamp 0
transform 1 0 26358 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_509
timestamp 0
transform 1 0 26450 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_511
timestamp 0
transform 1 0 26542 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_519
timestamp 0
transform 1 0 26910 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_527
timestamp 0
transform 1 0 27278 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_535
timestamp 0
transform 1 0 27646 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_543
timestamp 0
transform 1 0 28014 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_551
timestamp 0
transform 1 0 28382 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_88_559
timestamp 0
transform 1 0 28750 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_88_567
timestamp 0
transform 1 0 29118 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_569
timestamp 0
transform 1 0 29210 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_88_571
timestamp 0
transform 1 0 29302 0 1 27200
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_88_579
timestamp 0
transform 1 0 29670 0 1 27200
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_88_583
timestamp 0
transform 1 0 29854 0 1 27200
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_88_585
timestamp 0
transform 1 0 29946 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_89_0
timestamp 0
transform 1 0 3036 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_8
timestamp 0
transform 1 0 3404 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_16
timestamp 0
transform 1 0 3772 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_24
timestamp 0
transform 1 0 4140 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_56
timestamp 0
transform 1 0 5612 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_89_61
timestamp 0
transform 1 0 5842 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_69
timestamp 0
transform 1 0 6210 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_89_73
timestamp 0
transform 1 0 6394 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_89_77
timestamp 0
transform 1 0 6578 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_89_85
timestamp 0
transform 1 0 6946 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_89_95
timestamp 0
transform 1 0 7406 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_103
timestamp 0
transform 1 0 7774 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_111
timestamp 0
transform 1 0 8142 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_89_119
timestamp 0
transform 1 0 8510 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_89_121
timestamp 0
transform 1 0 8602 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_129
timestamp 0
transform 1 0 8970 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_137
timestamp 0
transform 1 0 9338 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_145
timestamp 0
transform 1 0 9706 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_153
timestamp 0
transform 1 0 10074 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_89_162
timestamp 0
transform 1 0 10488 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_170
timestamp 0
transform 1 0 10856 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_89_178
timestamp 0
transform 1 0 11224 0 -1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_89_181
timestamp 0
transform 1 0 11362 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_89_185
timestamp 0
transform 1 0 11546 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_89_189
timestamp 0
transform 1 0 11730 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_89_193
timestamp 0
transform 1 0 11914 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_89_203
timestamp 0
transform 1 0 12374 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_211
timestamp 0
transform 1 0 12742 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_219
timestamp 0
transform 1 0 13110 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 0
transform 1 0 13294 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_89_228
timestamp 0
transform 1 0 13524 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_236
timestamp 0
transform 1 0 13892 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_89_241
timestamp 0
transform 1 0 14122 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_249
timestamp 0
transform 1 0 14490 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_257
timestamp 0
transform 1 0 14858 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_89_261
timestamp 0
transform 1 0 15042 0 -1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_89_271
timestamp 0
transform 1 0 15502 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_89_278
timestamp 0
transform 1 0 15824 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_286
timestamp 0
transform 1 0 16192 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_294
timestamp 0
transform 1 0 16560 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_89_298
timestamp 0
transform 1 0 16744 0 -1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_89_301
timestamp 0
transform 1 0 16882 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_309
timestamp 0
transform 1 0 17250 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_317
timestamp 0
transform 1 0 17618 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_328
timestamp 0
transform 1 0 18124 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_89_341
timestamp 0
transform 1 0 18722 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_89_350
timestamp 0
transform 1 0 19136 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_89_358
timestamp 0
transform 1 0 19504 0 -1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_89_361
timestamp 0
transform 1 0 19642 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_369
timestamp 0
transform 1 0 20010 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_377
timestamp 0
transform 1 0 20378 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_385
timestamp 0
transform 1 0 20746 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_393
timestamp 0
transform 1 0 21114 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_401
timestamp 0
transform 1 0 21482 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_409
timestamp 0
transform 1 0 21850 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_89_417
timestamp 0
transform 1 0 22218 0 -1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_89_419
timestamp 0
transform 1 0 22310 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_89_421
timestamp 0
transform 1 0 22402 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_429
timestamp 0
transform 1 0 22770 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_437
timestamp 0
transform 1 0 23138 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_445
timestamp 0
transform 1 0 23506 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_453
timestamp 0
transform 1 0 23874 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_461
timestamp 0
transform 1 0 24242 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_469
timestamp 0
transform 1 0 24610 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_89_477
timestamp 0
transform 1 0 24978 0 -1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_89_479
timestamp 0
transform 1 0 25070 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_89_481
timestamp 0
transform 1 0 25162 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_489
timestamp 0
transform 1 0 25530 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_497
timestamp 0
transform 1 0 25898 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_505
timestamp 0
transform 1 0 26266 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_513
timestamp 0
transform 1 0 26634 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_521
timestamp 0
transform 1 0 27002 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_529
timestamp 0
transform 1 0 27370 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_89_537
timestamp 0
transform 1 0 27738 0 -1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_89_539
timestamp 0
transform 1 0 27830 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_89_541
timestamp 0
transform 1 0 27922 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_549
timestamp 0
transform 1 0 28290 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_557
timestamp 0
transform 1 0 28658 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_565
timestamp 0
transform 1 0 29026 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_89_573
timestamp 0
transform 1 0 29394 0 -1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_89_581
timestamp 0
transform 1 0 29762 0 -1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_89_585
timestamp 0
transform 1 0 29946 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_0
timestamp 0
transform 1 0 3036 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_8
timestamp 0
transform 1 0 3404 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_16
timestamp 0
transform 1 0 3772 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_90_24
timestamp 0
transform 1 0 4140 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_90_28
timestamp 0
transform 1 0 4324 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_90_31
timestamp 0
transform 1 0 4462 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_39
timestamp 0
transform 1 0 4830 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_47
timestamp 0
transform 1 0 5198 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_55
timestamp 0
transform 1 0 5566 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_63
timestamp 0
transform 1 0 5934 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_71
timestamp 0
transform 1 0 6302 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_79
timestamp 0
transform 1 0 6670 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_90_87
timestamp 0
transform 1 0 7038 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_89
timestamp 0
transform 1 0 7130 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_91
timestamp 0
transform 1 0 7222 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_99
timestamp 0
transform 1 0 7590 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_107
timestamp 0
transform 1 0 7958 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_115
timestamp 0
transform 1 0 8326 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_123
timestamp 0
transform 1 0 8694 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_131
timestamp 0
transform 1 0 9062 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_139
timestamp 0
transform 1 0 9430 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_90_147
timestamp 0
transform 1 0 9798 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_149
timestamp 0
transform 1 0 9890 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_151
timestamp 0
transform 1 0 9982 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_90_159
timestamp 0
transform 1 0 10350 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_163
timestamp 0
transform 1 0 10534 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_171
timestamp 0
transform 1 0 10902 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_90_179
timestamp 0
transform 1 0 11270 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_90_183
timestamp 0
transform 1 0 11454 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_185
timestamp 0
transform 1 0 11546 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_90_189
timestamp 0
transform 1 0 11730 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_90_204
timestamp 0
transform 1 0 12420 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_90_208
timestamp 0
transform 1 0 12604 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_90_211
timestamp 0
transform 1 0 12742 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_219
timestamp 0
transform 1 0 13110 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_227
timestamp 0
transform 1 0 13478 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_235
timestamp 0
transform 1 0 13846 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_243
timestamp 0
transform 1 0 14214 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_251
timestamp 0
transform 1 0 14582 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_259
timestamp 0
transform 1 0 14950 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_90_267
timestamp 0
transform 1 0 15318 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_269
timestamp 0
transform 1 0 15410 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_271
timestamp 0
transform 1 0 15502 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_279
timestamp 0
transform 1 0 15870 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_287
timestamp 0
transform 1 0 16238 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_295
timestamp 0
transform 1 0 16606 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_90_303
timestamp 0
transform 1 0 16974 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_90_314
timestamp 0
transform 1 0 17480 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_90_321
timestamp 0
transform 1 0 17802 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_90_329
timestamp 0
transform 1 0 18170 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_331
timestamp 0
transform 1 0 18262 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_90_339
timestamp 0
transform 1 0 18630 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_90_356
timestamp 0
transform 1 0 19412 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_90_363
timestamp 0
transform 1 0 19734 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_90_371
timestamp 0
transform 1 0 20102 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_90_375
timestamp 0
transform 1 0 20286 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_90_385
timestamp 0
transform 1 0 20746 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_90_389
timestamp 0
transform 1 0 20930 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_391
timestamp 0
transform 1 0 21022 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_399
timestamp 0
transform 1 0 21390 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_407
timestamp 0
transform 1 0 21758 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_415
timestamp 0
transform 1 0 22126 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_423
timestamp 0
transform 1 0 22494 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_431
timestamp 0
transform 1 0 22862 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_439
timestamp 0
transform 1 0 23230 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_90_447
timestamp 0
transform 1 0 23598 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_449
timestamp 0
transform 1 0 23690 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_451
timestamp 0
transform 1 0 23782 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_459
timestamp 0
transform 1 0 24150 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_467
timestamp 0
transform 1 0 24518 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_475
timestamp 0
transform 1 0 24886 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_483
timestamp 0
transform 1 0 25254 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_491
timestamp 0
transform 1 0 25622 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_499
timestamp 0
transform 1 0 25990 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_90_507
timestamp 0
transform 1 0 26358 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_509
timestamp 0
transform 1 0 26450 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_511
timestamp 0
transform 1 0 26542 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_519
timestamp 0
transform 1 0 26910 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_527
timestamp 0
transform 1 0 27278 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_535
timestamp 0
transform 1 0 27646 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_543
timestamp 0
transform 1 0 28014 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_551
timestamp 0
transform 1 0 28382 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_90_559
timestamp 0
transform 1 0 28750 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_90_567
timestamp 0
transform 1 0 29118 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_569
timestamp 0
transform 1 0 29210 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_90_571
timestamp 0
transform 1 0 29302 0 1 27744
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_90_579
timestamp 0
transform 1 0 29670 0 1 27744
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_90_583
timestamp 0
transform 1 0 29854 0 1 27744
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_90_585
timestamp 0
transform 1 0 29946 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_91_0
timestamp 0
transform 1 0 3036 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_8
timestamp 0
transform 1 0 3404 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_16
timestamp 0
transform 1 0 3772 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_24
timestamp 0
transform 1 0 4140 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_32
timestamp 0
transform 1 0 4508 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_91_40
timestamp 0
transform 1 0 4876 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_91_44
timestamp 0
transform 1 0 5060 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_91_46
timestamp 0
transform 1 0 5152 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_91_56
timestamp 0
transform 1 0 5612 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_91_61
timestamp 0
transform 1 0 5842 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_69
timestamp 0
transform 1 0 6210 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_77
timestamp 0
transform 1 0 6578 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_85
timestamp 0
transform 1 0 6946 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_93
timestamp 0
transform 1 0 7314 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_101
timestamp 0
transform 1 0 7682 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_109
timestamp 0
transform 1 0 8050 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_91_117
timestamp 0
transform 1 0 8418 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_91_119
timestamp 0
transform 1 0 8510 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_91_121
timestamp 0
transform 1 0 8602 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_91_131
timestamp 0
transform 1 0 9062 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_91_139
timestamp 0
transform 1 0 9430 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_91_143
timestamp 0
transform 1 0 9614 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_91_147
timestamp 0
transform 1 0 9798 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_91_151
timestamp 0
transform 1 0 9982 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_91_153
timestamp 0
transform 1 0 10074 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_91_158
timestamp 0
transform 1 0 10304 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_91_167
timestamp 0
transform 1 0 10718 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_91_175
timestamp 0
transform 1 0 11086 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_91_179
timestamp 0
transform 1 0 11270 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_91_181
timestamp 0
transform 1 0 11362 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_196
timestamp 0
transform 1 0 12052 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_204
timestamp 0
transform 1 0 12420 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_215
timestamp 0
transform 1 0 12926 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_226
timestamp 0
transform 1 0 13432 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_91_234
timestamp 0
transform 1 0 13800 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_91_238
timestamp 0
transform 1 0 13984 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_91_241
timestamp 0
transform 1 0 14122 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_91_253
timestamp 0
transform 1 0 14674 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_261
timestamp 0
transform 1 0 15042 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_279
timestamp 0
transform 1 0 15870 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_287
timestamp 0
transform 1 0 16238 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_91_295
timestamp 0
transform 1 0 16606 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_91_299
timestamp 0
transform 1 0 16790 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_91_301
timestamp 0
transform 1 0 16882 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_91_313
timestamp 0
transform 1 0 17434 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_91_323
timestamp 0
transform 1 0 17894 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_91_330
timestamp 0
transform 1 0 18216 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_91_338
timestamp 0
transform 1 0 18584 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_91_356
timestamp 0
transform 1 0 19412 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_91_361
timestamp 0
transform 1 0 19642 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_91_369
timestamp 0
transform 1 0 20010 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_91_393
timestamp 0
transform 1 0 21114 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_401
timestamp 0
transform 1 0 21482 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_409
timestamp 0
transform 1 0 21850 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_91_417
timestamp 0
transform 1 0 22218 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_91_419
timestamp 0
transform 1 0 22310 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_91_421
timestamp 0
transform 1 0 22402 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_429
timestamp 0
transform 1 0 22770 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_437
timestamp 0
transform 1 0 23138 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_445
timestamp 0
transform 1 0 23506 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_453
timestamp 0
transform 1 0 23874 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_461
timestamp 0
transform 1 0 24242 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_469
timestamp 0
transform 1 0 24610 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_91_477
timestamp 0
transform 1 0 24978 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_91_479
timestamp 0
transform 1 0 25070 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_91_481
timestamp 0
transform 1 0 25162 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_489
timestamp 0
transform 1 0 25530 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_497
timestamp 0
transform 1 0 25898 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_505
timestamp 0
transform 1 0 26266 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_513
timestamp 0
transform 1 0 26634 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_521
timestamp 0
transform 1 0 27002 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_529
timestamp 0
transform 1 0 27370 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_91_537
timestamp 0
transform 1 0 27738 0 -1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_91_539
timestamp 0
transform 1 0 27830 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_91_541
timestamp 0
transform 1 0 27922 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_549
timestamp 0
transform 1 0 28290 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_557
timestamp 0
transform 1 0 28658 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_565
timestamp 0
transform 1 0 29026 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_91_573
timestamp 0
transform 1 0 29394 0 -1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_91_581
timestamp 0
transform 1 0 29762 0 -1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_91_585
timestamp 0
transform 1 0 29946 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_92_0
timestamp 0
transform 1 0 3036 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_8
timestamp 0
transform 1 0 3404 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_16
timestamp 0
transform 1 0 3772 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_92_24
timestamp 0
transform 1 0 4140 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_92_28
timestamp 0
transform 1 0 4324 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_92_31
timestamp 0
transform 1 0 4462 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_92_39
timestamp 0
transform 1 0 4830 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_92_43
timestamp 0
transform 1 0 5014 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 0
transform 1 0 5106 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_92_55
timestamp 0
transform 1 0 5566 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_63
timestamp 0
transform 1 0 5934 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_71
timestamp 0
transform 1 0 6302 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_92_84
timestamp 0
transform 1 0 6900 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_92_88
timestamp 0
transform 1 0 7084 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_92_91
timestamp 0
transform 1 0 7222 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_99
timestamp 0
transform 1 0 7590 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_107
timestamp 0
transform 1 0 7958 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_92_115
timestamp 0
transform 1 0 8326 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_92_141
timestamp 0
transform 1 0 9522 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_92_149
timestamp 0
transform 1 0 9890 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_92_151
timestamp 0
transform 1 0 9982 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_92_171
timestamp 0
transform 1 0 10902 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_179
timestamp 0
transform 1 0 11270 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_187
timestamp 0
transform 1 0 11638 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_195
timestamp 0
transform 1 0 12006 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_92_203
timestamp 0
transform 1 0 12374 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_92_207
timestamp 0
transform 1 0 12558 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_92_209
timestamp 0
transform 1 0 12650 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_92_211
timestamp 0
transform 1 0 12742 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_92_238
timestamp 0
transform 1 0 13984 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_92_242
timestamp 0
transform 1 0 14168 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_92_266
timestamp 0
transform 1 0 15272 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_92_271
timestamp 0
transform 1 0 15502 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_92_284
timestamp 0
transform 1 0 16100 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_92_292
timestamp 0
transform 1 0 16468 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_92_294
timestamp 0
transform 1 0 16560 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_92_304
timestamp 0
transform 1 0 17020 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_92_324
timestamp 0
transform 1 0 17940 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_92_328
timestamp 0
transform 1 0 18124 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_92_331
timestamp 0
transform 1 0 18262 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_339
timestamp 0
transform 1 0 18630 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_92_347
timestamp 0
transform 1 0 18998 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_92_351
timestamp 0
transform 1 0 19182 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_92_363
timestamp 0
transform 1 0 19734 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_92_371
timestamp 0
transform 1 0 20102 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_92_384
timestamp 0
transform 1 0 20700 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_92_388
timestamp 0
transform 1 0 20884 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_92_391
timestamp 0
transform 1 0 21022 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_399
timestamp 0
transform 1 0 21390 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_407
timestamp 0
transform 1 0 21758 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_415
timestamp 0
transform 1 0 22126 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_423
timestamp 0
transform 1 0 22494 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_431
timestamp 0
transform 1 0 22862 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_439
timestamp 0
transform 1 0 23230 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_92_447
timestamp 0
transform 1 0 23598 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_92_449
timestamp 0
transform 1 0 23690 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_92_451
timestamp 0
transform 1 0 23782 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_459
timestamp 0
transform 1 0 24150 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_467
timestamp 0
transform 1 0 24518 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_475
timestamp 0
transform 1 0 24886 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_483
timestamp 0
transform 1 0 25254 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_491
timestamp 0
transform 1 0 25622 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_499
timestamp 0
transform 1 0 25990 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_92_507
timestamp 0
transform 1 0 26358 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_92_509
timestamp 0
transform 1 0 26450 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_92_511
timestamp 0
transform 1 0 26542 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_519
timestamp 0
transform 1 0 26910 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_527
timestamp 0
transform 1 0 27278 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_535
timestamp 0
transform 1 0 27646 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_543
timestamp 0
transform 1 0 28014 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_551
timestamp 0
transform 1 0 28382 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_92_559
timestamp 0
transform 1 0 28750 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_92_567
timestamp 0
transform 1 0 29118 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_92_569
timestamp 0
transform 1 0 29210 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_92_571
timestamp 0
transform 1 0 29302 0 1 28288
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_92_579
timestamp 0
transform 1 0 29670 0 1 28288
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_92_583
timestamp 0
transform 1 0 29854 0 1 28288
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_92_585
timestamp 0
transform 1 0 29946 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_93_0
timestamp 0
transform 1 0 3036 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_8
timestamp 0
transform 1 0 3404 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_16
timestamp 0
transform 1 0 3772 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_24
timestamp 0
transform 1 0 4140 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_32
timestamp 0
transform 1 0 4508 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_93_56
timestamp 0
transform 1 0 5612 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_93_61
timestamp 0
transform 1 0 5842 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_93_69
timestamp 0
transform 1 0 6210 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_93_79
timestamp 0
transform 1 0 6670 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_93_87
timestamp 0
transform 1 0 7038 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_95
timestamp 0
transform 1 0 7406 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_103
timestamp 0
transform 1 0 7774 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_93_107
timestamp 0
transform 1 0 7958 0 -1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_93_109
timestamp 0
transform 1 0 8050 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_93_116
timestamp 0
transform 1 0 8372 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_93_121
timestamp 0
transform 1 0 8602 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_93_128
timestamp 0
transform 1 0 8924 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_136
timestamp 0
transform 1 0 9292 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_144
timestamp 0
transform 1 0 9660 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_152
timestamp 0
transform 1 0 10028 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_93_156
timestamp 0
transform 1 0 10212 0 -1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_93_162
timestamp 0
transform 1 0 10488 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_170
timestamp 0
transform 1 0 10856 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_93_178
timestamp 0
transform 1 0 11224 0 -1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_93_181
timestamp 0
transform 1 0 11362 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_189
timestamp 0
transform 1 0 11730 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_197
timestamp 0
transform 1 0 12098 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_205
timestamp 0
transform 1 0 12466 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_213
timestamp 0
transform 1 0 12834 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_93_221
timestamp 0
transform 1 0 13202 0 -1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 0
transform 1 0 13294 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_93_228
timestamp 0
transform 1 0 13524 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_236
timestamp 0
transform 1 0 13892 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_93_241
timestamp 0
transform 1 0 14122 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_249
timestamp 0
transform 1 0 14490 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_257
timestamp 0
transform 1 0 14858 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_265
timestamp 0
transform 1 0 15226 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_273
timestamp 0
transform 1 0 15594 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_93_280
timestamp 0
transform 1 0 15916 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_288
timestamp 0
transform 1 0 16284 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_296
timestamp 0
transform 1 0 16652 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_93_301
timestamp 0
transform 1 0 16882 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_93_309
timestamp 0
transform 1 0 17250 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_93_336
timestamp 0
transform 1 0 18492 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_344
timestamp 0
transform 1 0 18860 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_352
timestamp 0
transform 1 0 19228 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_361
timestamp 0
transform 1 0 19642 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_93_369
timestamp 0
transform 1 0 20010 0 -1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_93_371
timestamp 0
transform 1 0 20102 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_93_392
timestamp 0
transform 1 0 21068 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_400
timestamp 0
transform 1 0 21436 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_408
timestamp 0
transform 1 0 21804 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_416
timestamp 0
transform 1 0 22172 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_93_421
timestamp 0
transform 1 0 22402 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_429
timestamp 0
transform 1 0 22770 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_437
timestamp 0
transform 1 0 23138 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_445
timestamp 0
transform 1 0 23506 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_453
timestamp 0
transform 1 0 23874 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_461
timestamp 0
transform 1 0 24242 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_469
timestamp 0
transform 1 0 24610 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_93_477
timestamp 0
transform 1 0 24978 0 -1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_93_479
timestamp 0
transform 1 0 25070 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_93_481
timestamp 0
transform 1 0 25162 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_489
timestamp 0
transform 1 0 25530 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_497
timestamp 0
transform 1 0 25898 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_505
timestamp 0
transform 1 0 26266 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_513
timestamp 0
transform 1 0 26634 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_521
timestamp 0
transform 1 0 27002 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_529
timestamp 0
transform 1 0 27370 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_93_537
timestamp 0
transform 1 0 27738 0 -1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_93_539
timestamp 0
transform 1 0 27830 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_93_541
timestamp 0
transform 1 0 27922 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_549
timestamp 0
transform 1 0 28290 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_557
timestamp 0
transform 1 0 28658 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_565
timestamp 0
transform 1 0 29026 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_93_573
timestamp 0
transform 1 0 29394 0 -1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_93_581
timestamp 0
transform 1 0 29762 0 -1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_93_585
timestamp 0
transform 1 0 29946 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_0
timestamp 0
transform 1 0 3036 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_8
timestamp 0
transform 1 0 3404 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_16
timestamp 0
transform 1 0 3772 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_24
timestamp 0
transform 1 0 4140 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_28
timestamp 0
transform 1 0 4324 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_94_31
timestamp 0
transform 1 0 4462 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_35
timestamp 0
transform 1 0 4646 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_37
timestamp 0
transform 1 0 4738 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_58
timestamp 0
transform 1 0 5704 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_66
timestamp 0
transform 1 0 6072 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_74
timestamp 0
transform 1 0 6440 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_78
timestamp 0
transform 1 0 6624 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_94_86
timestamp 0
transform 1 0 6992 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_94_91
timestamp 0
transform 1 0 7222 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_94_98
timestamp 0
transform 1 0 7544 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_106
timestamp 0
transform 1 0 7912 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_94_114
timestamp 0
transform 1 0 8280 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_116
timestamp 0
transform 1 0 8372 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_94_120
timestamp 0
transform 1 0 8556 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_94_130
timestamp 0
transform 1 0 9016 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_138
timestamp 0
transform 1 0 9384 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_146
timestamp 0
transform 1 0 9752 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_94_151
timestamp 0
transform 1 0 9982 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_155
timestamp 0
transform 1 0 10166 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_94_161
timestamp 0
transform 1 0 10442 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_169
timestamp 0
transform 1 0 10810 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_173
timestamp 0
transform 1 0 10994 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_94_182
timestamp 0
transform 1 0 11408 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_186
timestamp 0
transform 1 0 11592 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_94_193
timestamp 0
transform 1 0 11914 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_201
timestamp 0
transform 1 0 12282 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_94_209
timestamp 0
transform 1 0 12650 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_211
timestamp 0
transform 1 0 12742 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_219
timestamp 0
transform 1 0 13110 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_227
timestamp 0
transform 1 0 13478 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_231
timestamp 0
transform 1 0 13662 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_94_236
timestamp 0
transform 1 0 13892 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_94_243
timestamp 0
transform 1 0 14214 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_251
timestamp 0
transform 1 0 14582 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_259
timestamp 0
transform 1 0 14950 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_94_266
timestamp 0
transform 1 0 15272 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_94_271
timestamp 0
transform 1 0 15502 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_94_279
timestamp 0
transform 1 0 15870 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_283
timestamp 0
transform 1 0 16054 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_285
timestamp 0
transform 1 0 16146 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_291
timestamp 0
transform 1 0 16422 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_299
timestamp 0
transform 1 0 16790 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_94_309
timestamp 0
transform 1 0 17250 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_94_318
timestamp 0
transform 1 0 17664 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_326
timestamp 0
transform 1 0 18032 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_94_331
timestamp 0
transform 1 0 18262 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_339
timestamp 0
transform 1 0 18630 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_347
timestamp 0
transform 1 0 18998 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_355
timestamp 0
transform 1 0 19366 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_363
timestamp 0
transform 1 0 19734 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_371
timestamp 0
transform 1 0 20102 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_379
timestamp 0
transform 1 0 20470 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_94_387
timestamp 0
transform 1 0 20838 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_389
timestamp 0
transform 1 0 20930 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_391
timestamp 0
transform 1 0 21022 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_399
timestamp 0
transform 1 0 21390 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_407
timestamp 0
transform 1 0 21758 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_415
timestamp 0
transform 1 0 22126 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_423
timestamp 0
transform 1 0 22494 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_431
timestamp 0
transform 1 0 22862 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_439
timestamp 0
transform 1 0 23230 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_94_447
timestamp 0
transform 1 0 23598 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_449
timestamp 0
transform 1 0 23690 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_451
timestamp 0
transform 1 0 23782 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_459
timestamp 0
transform 1 0 24150 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_467
timestamp 0
transform 1 0 24518 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_475
timestamp 0
transform 1 0 24886 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_483
timestamp 0
transform 1 0 25254 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_491
timestamp 0
transform 1 0 25622 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_499
timestamp 0
transform 1 0 25990 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_94_507
timestamp 0
transform 1 0 26358 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_509
timestamp 0
transform 1 0 26450 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_511
timestamp 0
transform 1 0 26542 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_519
timestamp 0
transform 1 0 26910 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_527
timestamp 0
transform 1 0 27278 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_535
timestamp 0
transform 1 0 27646 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_543
timestamp 0
transform 1 0 28014 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_551
timestamp 0
transform 1 0 28382 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_94_559
timestamp 0
transform 1 0 28750 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_94_567
timestamp 0
transform 1 0 29118 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_569
timestamp 0
transform 1 0 29210 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_94_571
timestamp 0
transform 1 0 29302 0 1 28832
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_94_579
timestamp 0
transform 1 0 29670 0 1 28832
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_94_583
timestamp 0
transform 1 0 29854 0 1 28832
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_94_585
timestamp 0
transform 1 0 29946 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_95_0
timestamp 0
transform 1 0 3036 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_8
timestamp 0
transform 1 0 3404 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_16
timestamp 0
transform 1 0 3772 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_24
timestamp 0
transform 1 0 4140 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_32
timestamp 0
transform 1 0 4508 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_40
timestamp 0
transform 1 0 4876 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_48
timestamp 0
transform 1 0 5244 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_95_56
timestamp 0
transform 1 0 5612 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_95_61
timestamp 0
transform 1 0 5842 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_69
timestamp 0
transform 1 0 6210 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_95_77
timestamp 0
transform 1 0 6578 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_95_81
timestamp 0
transform 1 0 6762 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_95_106
timestamp 0
transform 1 0 7912 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_95_114
timestamp 0
transform 1 0 8280 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_95_118
timestamp 0
transform 1 0 8464 0 -1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_4  FILLER_95_121
timestamp 0
transform 1 0 8602 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_95_125
timestamp 0
transform 1 0 8786 0 -1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_95_130
timestamp 0
transform 1 0 9016 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_138
timestamp 0
transform 1 0 9384 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_95_146
timestamp 0
transform 1 0 9752 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_95_150
timestamp 0
transform 1 0 9936 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_95_167
timestamp 0
transform 1 0 10718 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_95_175
timestamp 0
transform 1 0 11086 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_95_179
timestamp 0
transform 1 0 11270 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_95_181
timestamp 0
transform 1 0 11362 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_95_185
timestamp 0
transform 1 0 11546 0 -1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_95_203
timestamp 0
transform 1 0 12374 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_211
timestamp 0
transform 1 0 12742 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_95_219
timestamp 0
transform 1 0 13110 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_95_236
timestamp 0
transform 1 0 13892 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_95_241
timestamp 0
transform 1 0 14122 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_95_249
timestamp 0
transform 1 0 14490 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_95_255
timestamp 0
transform 1 0 14766 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_95_259
timestamp 0
transform 1 0 14950 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_95_276
timestamp 0
transform 1 0 15732 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_95_296
timestamp 0
transform 1 0 16652 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_95_301
timestamp 0
transform 1 0 16882 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_309
timestamp 0
transform 1 0 17250 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_317
timestamp 0
transform 1 0 17618 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_325
timestamp 0
transform 1 0 17986 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_333
timestamp 0
transform 1 0 18354 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_341
timestamp 0
transform 1 0 18722 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_349
timestamp 0
transform 1 0 19090 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_95_357
timestamp 0
transform 1 0 19458 0 -1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_95_359
timestamp 0
transform 1 0 19550 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_95_361
timestamp 0
transform 1 0 19642 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_369
timestamp 0
transform 1 0 20010 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_377
timestamp 0
transform 1 0 20378 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_385
timestamp 0
transform 1 0 20746 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_393
timestamp 0
transform 1 0 21114 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_401
timestamp 0
transform 1 0 21482 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_409
timestamp 0
transform 1 0 21850 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_95_417
timestamp 0
transform 1 0 22218 0 -1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_95_419
timestamp 0
transform 1 0 22310 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_95_421
timestamp 0
transform 1 0 22402 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_429
timestamp 0
transform 1 0 22770 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_437
timestamp 0
transform 1 0 23138 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_445
timestamp 0
transform 1 0 23506 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_453
timestamp 0
transform 1 0 23874 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_461
timestamp 0
transform 1 0 24242 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_469
timestamp 0
transform 1 0 24610 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_95_477
timestamp 0
transform 1 0 24978 0 -1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_95_479
timestamp 0
transform 1 0 25070 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_95_481
timestamp 0
transform 1 0 25162 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_489
timestamp 0
transform 1 0 25530 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_497
timestamp 0
transform 1 0 25898 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_505
timestamp 0
transform 1 0 26266 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_513
timestamp 0
transform 1 0 26634 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_521
timestamp 0
transform 1 0 27002 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_529
timestamp 0
transform 1 0 27370 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_95_537
timestamp 0
transform 1 0 27738 0 -1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_95_539
timestamp 0
transform 1 0 27830 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_95_541
timestamp 0
transform 1 0 27922 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_549
timestamp 0
transform 1 0 28290 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_557
timestamp 0
transform 1 0 28658 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_565
timestamp 0
transform 1 0 29026 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_95_573
timestamp 0
transform 1 0 29394 0 -1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_95_581
timestamp 0
transform 1 0 29762 0 -1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_95_585
timestamp 0
transform 1 0 29946 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_0
timestamp 0
transform 1 0 3036 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_8
timestamp 0
transform 1 0 3404 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_16
timestamp 0
transform 1 0 3772 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_96_24
timestamp 0
transform 1 0 4140 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_96_28
timestamp 0
transform 1 0 4324 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_96_31
timestamp 0
transform 1 0 4462 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_39
timestamp 0
transform 1 0 4830 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_47
timestamp 0
transform 1 0 5198 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_55
timestamp 0
transform 1 0 5566 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_63
timestamp 0
transform 1 0 5934 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_71
timestamp 0
transform 1 0 6302 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_79
timestamp 0
transform 1 0 6670 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_87
timestamp 0
transform 1 0 7038 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_89
timestamp 0
transform 1 0 7130 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_91
timestamp 0
transform 1 0 7222 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_99
timestamp 0
transform 1 0 7590 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_107
timestamp 0
transform 1 0 7958 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_115
timestamp 0
transform 1 0 8326 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_123
timestamp 0
transform 1 0 8694 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_131
timestamp 0
transform 1 0 9062 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_139
timestamp 0
transform 1 0 9430 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_147
timestamp 0
transform 1 0 9798 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_149
timestamp 0
transform 1 0 9890 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_96_151
timestamp 0
transform 1 0 9982 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_96_155
timestamp 0
transform 1 0 10166 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_96_161
timestamp 0
transform 1 0 10442 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_169
timestamp 0
transform 1 0 10810 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_177
timestamp 0
transform 1 0 11178 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_185
timestamp 0
transform 1 0 11546 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_187
timestamp 0
transform 1 0 11638 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_96_192
timestamp 0
transform 1 0 11868 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_8  FILLER_96_199
timestamp 0
transform 1 0 12190 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_207
timestamp 0
transform 1 0 12558 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_209
timestamp 0
transform 1 0 12650 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_211
timestamp 0
transform 1 0 12742 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_219
timestamp 0
transform 1 0 13110 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_227
timestamp 0
transform 1 0 13478 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_235
timestamp 0
transform 1 0 13846 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_243
timestamp 0
transform 1 0 14214 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_251
timestamp 0
transform 1 0 14582 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_259
timestamp 0
transform 1 0 14950 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_267
timestamp 0
transform 1 0 15318 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_269
timestamp 0
transform 1 0 15410 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_4  FILLER_96_271
timestamp 0
transform 1 0 15502 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_4  FILLER_96_279
timestamp 0
transform 1 0 15870 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_96_283
timestamp 0
transform 1 0 16054 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_288
timestamp 0
transform 1 0 16284 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_296
timestamp 0
transform 1 0 16652 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_304
timestamp 0
transform 1 0 17020 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_312
timestamp 0
transform 1 0 17388 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_320
timestamp 0
transform 1 0 17756 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_328
timestamp 0
transform 1 0 18124 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_96_331
timestamp 0
transform 1 0 18262 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_339
timestamp 0
transform 1 0 18630 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_347
timestamp 0
transform 1 0 18998 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_355
timestamp 0
transform 1 0 19366 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_363
timestamp 0
transform 1 0 19734 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_371
timestamp 0
transform 1 0 20102 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_379
timestamp 0
transform 1 0 20470 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_387
timestamp 0
transform 1 0 20838 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_389
timestamp 0
transform 1 0 20930 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_391
timestamp 0
transform 1 0 21022 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_399
timestamp 0
transform 1 0 21390 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_407
timestamp 0
transform 1 0 21758 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_415
timestamp 0
transform 1 0 22126 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_423
timestamp 0
transform 1 0 22494 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_431
timestamp 0
transform 1 0 22862 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_439
timestamp 0
transform 1 0 23230 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_447
timestamp 0
transform 1 0 23598 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_449
timestamp 0
transform 1 0 23690 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_451
timestamp 0
transform 1 0 23782 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_459
timestamp 0
transform 1 0 24150 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_467
timestamp 0
transform 1 0 24518 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_475
timestamp 0
transform 1 0 24886 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_483
timestamp 0
transform 1 0 25254 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_491
timestamp 0
transform 1 0 25622 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_499
timestamp 0
transform 1 0 25990 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_507
timestamp 0
transform 1 0 26358 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_509
timestamp 0
transform 1 0 26450 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_511
timestamp 0
transform 1 0 26542 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_519
timestamp 0
transform 1 0 26910 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_527
timestamp 0
transform 1 0 27278 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_535
timestamp 0
transform 1 0 27646 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_543
timestamp 0
transform 1 0 28014 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_551
timestamp 0
transform 1 0 28382 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_96_559
timestamp 0
transform 1 0 28750 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_2  FILLER_96_567
timestamp 0
transform 1 0 29118 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_569
timestamp 0
transform 1 0 29210 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_96_571
timestamp 0
transform 1 0 29302 0 1 29376
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_96_579
timestamp 0
transform 1 0 29670 0 1 29376
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_96_583
timestamp 0
transform 1 0 29854 0 1 29376
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_96_585
timestamp 0
transform 1 0 29946 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_0
timestamp 0
transform 1 0 3036 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_8
timestamp 0
transform 1 0 3404 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_16
timestamp 0
transform 1 0 3772 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_24
timestamp 0
transform 1 0 4140 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_97_28
timestamp 0
transform 1 0 4324 0 -1 29920
box 0 -24 92 296
use sky130_fd_sc_hd__fill_8  FILLER_97_31
timestamp 0
transform 1 0 4462 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_39
timestamp 0
transform 1 0 4830 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_47
timestamp 0
transform 1 0 5198 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_55
timestamp 0
transform 1 0 5566 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_59
timestamp 0
transform 1 0 5750 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_61
timestamp 0
transform 1 0 5842 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_69
timestamp 0
transform 1 0 6210 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_77
timestamp 0
transform 1 0 6578 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_85
timestamp 0
transform 1 0 6946 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_89
timestamp 0
transform 1 0 7130 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_91
timestamp 0
transform 1 0 7222 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_99
timestamp 0
transform 1 0 7590 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_107
timestamp 0
transform 1 0 7958 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_115
timestamp 0
transform 1 0 8326 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_119
timestamp 0
transform 1 0 8510 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_121
timestamp 0
transform 1 0 8602 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_129
timestamp 0
transform 1 0 8970 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_137
timestamp 0
transform 1 0 9338 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_145
timestamp 0
transform 1 0 9706 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_149
timestamp 0
transform 1 0 9890 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_151
timestamp 0
transform 1 0 9982 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_159
timestamp 0
transform 1 0 10350 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_167
timestamp 0
transform 1 0 10718 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_175
timestamp 0
transform 1 0 11086 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_179
timestamp 0
transform 1 0 11270 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_181
timestamp 0
transform 1 0 11362 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_189
timestamp 0
transform 1 0 11730 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_197
timestamp 0
transform 1 0 12098 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_205
timestamp 0
transform 1 0 12466 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_209
timestamp 0
transform 1 0 12650 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_211
timestamp 0
transform 1 0 12742 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_219
timestamp 0
transform 1 0 13110 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_227
timestamp 0
transform 1 0 13478 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_235
timestamp 0
transform 1 0 13846 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_239
timestamp 0
transform 1 0 14030 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_241
timestamp 0
transform 1 0 14122 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_249
timestamp 0
transform 1 0 14490 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_257
timestamp 0
transform 1 0 14858 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_265
timestamp 0
transform 1 0 15226 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_269
timestamp 0
transform 1 0 15410 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_271
timestamp 0
transform 1 0 15502 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 0
transform 1 0 15870 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_283
timestamp 0
transform 1 0 16054 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_291
timestamp 0
transform 1 0 16422 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_1  FILLER_97_299
timestamp 0
transform 1 0 16790 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_301
timestamp 0
transform 1 0 16882 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_309
timestamp 0
transform 1 0 17250 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_317
timestamp 0
transform 1 0 17618 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_325
timestamp 0
transform 1 0 17986 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_329
timestamp 0
transform 1 0 18170 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_331
timestamp 0
transform 1 0 18262 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_339
timestamp 0
transform 1 0 18630 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_347
timestamp 0
transform 1 0 18998 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_355
timestamp 0
transform 1 0 19366 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_359
timestamp 0
transform 1 0 19550 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_361
timestamp 0
transform 1 0 19642 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_369
timestamp 0
transform 1 0 20010 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_377
timestamp 0
transform 1 0 20378 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_385
timestamp 0
transform 1 0 20746 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_389
timestamp 0
transform 1 0 20930 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_391
timestamp 0
transform 1 0 21022 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_399
timestamp 0
transform 1 0 21390 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_407
timestamp 0
transform 1 0 21758 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_415
timestamp 0
transform 1 0 22126 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_419
timestamp 0
transform 1 0 22310 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_421
timestamp 0
transform 1 0 22402 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_429
timestamp 0
transform 1 0 22770 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_437
timestamp 0
transform 1 0 23138 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_445
timestamp 0
transform 1 0 23506 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_449
timestamp 0
transform 1 0 23690 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_451
timestamp 0
transform 1 0 23782 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_459
timestamp 0
transform 1 0 24150 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_467
timestamp 0
transform 1 0 24518 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_475
timestamp 0
transform 1 0 24886 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_479
timestamp 0
transform 1 0 25070 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_481
timestamp 0
transform 1 0 25162 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_489
timestamp 0
transform 1 0 25530 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_497
timestamp 0
transform 1 0 25898 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_505
timestamp 0
transform 1 0 26266 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_509
timestamp 0
transform 1 0 26450 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_511
timestamp 0
transform 1 0 26542 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_519
timestamp 0
transform 1 0 26910 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_527
timestamp 0
transform 1 0 27278 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_535
timestamp 0
transform 1 0 27646 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_539
timestamp 0
transform 1 0 27830 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_541
timestamp 0
transform 1 0 27922 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_549
timestamp 0
transform 1 0 28290 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_8  FILLER_97_557
timestamp 0
transform 1 0 28658 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_565
timestamp 0
transform 1 0 29026 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_1  FILLER_97_569
timestamp 0
transform 1 0 29210 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__fill_8  FILLER_97_571
timestamp 0
transform 1 0 29302 0 -1 29920
box 0 -24 368 296
use sky130_fd_sc_hd__fill_4  FILLER_97_579
timestamp 0
transform 1 0 29670 0 -1 29920
box 0 -24 184 296
use sky130_fd_sc_hd__fill_2  FILLER_97_583
timestamp 0
transform 1 0 29854 0 -1 29920
box 0 -24 92 296
use sky130_fd_sc_hd__fill_1  FILLER_97_585
timestamp 0
transform 1 0 29946 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__clkbuf_4  load_slew2
timestamp 0
transform 1 0 15686 0 1 24480
box 0 -24 276 296
use sky130_fd_sc_hd__buf_12  load_slew3
timestamp 0
transform 1 0 7406 0 1 16320
box 0 -24 736 296
use sky130_fd_sc_hd__buf_12  load_slew4
timestamp 0
transform 1 0 11868 0 -1 11968
box 0 -24 736 296
use sky130_fd_sc_hd__buf_16  load_slew5
timestamp 0
transform 1 0 10074 0 -1 12512
box 0 -24 1012 296
use sky130_fd_sc_hd__buf_16  load_slew6
timestamp 0
transform 1 0 6072 0 -1 11968
box 0 -24 1012 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_0
timestamp 0
transform 1 0 4416 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_1
timestamp 0
transform 1 0 5796 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_2
timestamp 0
transform 1 0 7176 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_3
timestamp 0
transform 1 0 8556 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_4
timestamp 0
transform 1 0 9936 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_5
timestamp 0
transform 1 0 11316 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_6
timestamp 0
transform 1 0 12696 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_7
timestamp 0
transform 1 0 14076 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_8
timestamp 0
transform 1 0 15456 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_9
timestamp 0
transform 1 0 16836 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_10
timestamp 0
transform 1 0 18216 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_11
timestamp 0
transform 1 0 19596 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_12
timestamp 0
transform 1 0 20976 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_13
timestamp 0
transform 1 0 22356 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_14
timestamp 0
transform 1 0 23736 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_15
timestamp 0
transform 1 0 25116 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_16
timestamp 0
transform 1 0 26496 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_17
timestamp 0
transform 1 0 27876 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_18
timestamp 0
transform 1 0 29256 0 1 3264
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_19
timestamp 0
transform 1 0 5796 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_20
timestamp 0
transform 1 0 8556 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_21
timestamp 0
transform 1 0 11316 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 0
transform 1 0 14076 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_23
timestamp 0
transform 1 0 16836 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_24
timestamp 0
transform 1 0 19596 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_25
timestamp 0
transform 1 0 22356 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_26
timestamp 0
transform 1 0 25116 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_27
timestamp 0
transform 1 0 27876 0 -1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_28
timestamp 0
transform 1 0 4416 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp 0
transform 1 0 7176 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_30
timestamp 0
transform 1 0 9936 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp 0
transform 1 0 12696 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_32
timestamp 0
transform 1 0 15456 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_33
timestamp 0
transform 1 0 18216 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_34
timestamp 0
transform 1 0 20976 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_35
timestamp 0
transform 1 0 23736 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_36
timestamp 0
transform 1 0 26496 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_37
timestamp 0
transform 1 0 29256 0 1 3808
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_38
timestamp 0
transform 1 0 5796 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_39
timestamp 0
transform 1 0 8556 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 0
transform 1 0 11316 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_41
timestamp 0
transform 1 0 14076 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp 0
transform 1 0 16836 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_43
timestamp 0
transform 1 0 19596 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_44
timestamp 0
transform 1 0 22356 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_45
timestamp 0
transform 1 0 25116 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_46
timestamp 0
transform 1 0 27876 0 -1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_47
timestamp 0
transform 1 0 4416 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_48
timestamp 0
transform 1 0 7176 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_49
timestamp 0
transform 1 0 9936 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_50
timestamp 0
transform 1 0 12696 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_51
timestamp 0
transform 1 0 15456 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_52
timestamp 0
transform 1 0 18216 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_53
timestamp 0
transform 1 0 20976 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_54
timestamp 0
transform 1 0 23736 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp 0
transform 1 0 26496 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp 0
transform 1 0 29256 0 1 4352
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_57
timestamp 0
transform 1 0 5796 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_58
timestamp 0
transform 1 0 8556 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_59
timestamp 0
transform 1 0 11316 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_60
timestamp 0
transform 1 0 14076 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_61
timestamp 0
transform 1 0 16836 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_62
timestamp 0
transform 1 0 19596 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_63
timestamp 0
transform 1 0 22356 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_64
timestamp 0
transform 1 0 25116 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp 0
transform 1 0 27876 0 -1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_66
timestamp 0
transform 1 0 4416 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp 0
transform 1 0 7176 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp 0
transform 1 0 9936 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp 0
transform 1 0 12696 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_70
timestamp 0
transform 1 0 15456 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp 0
transform 1 0 18216 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_72
timestamp 0
transform 1 0 20976 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp 0
transform 1 0 23736 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp 0
transform 1 0 26496 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp 0
transform 1 0 29256 0 1 4896
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp 0
transform 1 0 5796 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp 0
transform 1 0 8556 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_78
timestamp 0
transform 1 0 11316 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_79
timestamp 0
transform 1 0 14076 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 0
transform 1 0 16836 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 0
transform 1 0 19596 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 0
transform 1 0 22356 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp 0
transform 1 0 25116 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp 0
transform 1 0 27876 0 -1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 0
transform 1 0 4416 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_86
timestamp 0
transform 1 0 7176 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp 0
transform 1 0 9936 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp 0
transform 1 0 12696 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 0
transform 1 0 15456 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 0
transform 1 0 18216 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 0
transform 1 0 20976 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp 0
transform 1 0 23736 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp 0
transform 1 0 26496 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_94
timestamp 0
transform 1 0 29256 0 1 5440
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp 0
transform 1 0 5796 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp 0
transform 1 0 8556 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp 0
transform 1 0 11316 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp 0
transform 1 0 14076 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp 0
transform 1 0 16836 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp 0
transform 1 0 19596 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_101
timestamp 0
transform 1 0 22356 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_102
timestamp 0
transform 1 0 25116 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp 0
transform 1 0 27876 0 -1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp 0
transform 1 0 4416 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp 0
transform 1 0 7176 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp 0
transform 1 0 9936 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp 0
transform 1 0 12696 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp 0
transform 1 0 15456 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp 0
transform 1 0 18216 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_110
timestamp 0
transform 1 0 20976 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_111
timestamp 0
transform 1 0 23736 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp 0
transform 1 0 26496 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp 0
transform 1 0 29256 0 1 5984
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp 0
transform 1 0 5796 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp 0
transform 1 0 8556 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp 0
transform 1 0 11316 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp 0
transform 1 0 14076 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp 0
transform 1 0 16836 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp 0
transform 1 0 19596 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp 0
transform 1 0 22356 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp 0
transform 1 0 25116 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp 0
transform 1 0 27876 0 -1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_123
timestamp 0
transform 1 0 4416 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_124
timestamp 0
transform 1 0 7176 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_125
timestamp 0
transform 1 0 9936 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_126
timestamp 0
transform 1 0 12696 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_127
timestamp 0
transform 1 0 15456 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_128
timestamp 0
transform 1 0 18216 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_129
timestamp 0
transform 1 0 20976 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_130
timestamp 0
transform 1 0 23736 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_131
timestamp 0
transform 1 0 26496 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_132
timestamp 0
transform 1 0 29256 0 1 6528
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_133
timestamp 0
transform 1 0 5796 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_134
timestamp 0
transform 1 0 8556 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_135
timestamp 0
transform 1 0 11316 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_136
timestamp 0
transform 1 0 14076 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_137
timestamp 0
transform 1 0 16836 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_138
timestamp 0
transform 1 0 19596 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_139
timestamp 0
transform 1 0 22356 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 0
transform 1 0 25116 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 0
transform 1 0 27876 0 -1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_142
timestamp 0
transform 1 0 4416 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_143
timestamp 0
transform 1 0 7176 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 0
transform 1 0 9936 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 0
transform 1 0 12696 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 0
transform 1 0 15456 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 0
transform 1 0 18216 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_148
timestamp 0
transform 1 0 20976 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_149
timestamp 0
transform 1 0 23736 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 0
transform 1 0 26496 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 0
transform 1 0 29256 0 1 7072
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_152
timestamp 0
transform 1 0 5796 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_153
timestamp 0
transform 1 0 8556 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_154
timestamp 0
transform 1 0 11316 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_155
timestamp 0
transform 1 0 14076 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 0
transform 1 0 16836 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 0
transform 1 0 19596 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 0
transform 1 0 22356 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 0
transform 1 0 25116 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 0
transform 1 0 27876 0 -1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 0
transform 1 0 4416 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 0
transform 1 0 7176 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 0
transform 1 0 9936 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 0
transform 1 0 12696 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 0
transform 1 0 15456 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 0
transform 1 0 18216 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_167
timestamp 0
transform 1 0 20976 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_168
timestamp 0
transform 1 0 23736 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_169
timestamp 0
transform 1 0 26496 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_170
timestamp 0
transform 1 0 29256 0 1 7616
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 0
transform 1 0 5796 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_172
timestamp 0
transform 1 0 8556 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_173
timestamp 0
transform 1 0 11316 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_174
timestamp 0
transform 1 0 14076 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_175
timestamp 0
transform 1 0 16836 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_176
timestamp 0
transform 1 0 19596 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 0
transform 1 0 22356 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 0
transform 1 0 25116 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 0
transform 1 0 27876 0 -1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_180
timestamp 0
transform 1 0 4416 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_181
timestamp 0
transform 1 0 7176 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 0
transform 1 0 9936 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 0
transform 1 0 12696 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 0
transform 1 0 15456 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 0
transform 1 0 18216 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 0
transform 1 0 20976 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 0
transform 1 0 23736 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_188
timestamp 0
transform 1 0 26496 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_189
timestamp 0
transform 1 0 29256 0 1 8160
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 0
transform 1 0 5796 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 0
transform 1 0 8556 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 0
transform 1 0 11316 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_193
timestamp 0
transform 1 0 14076 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_194
timestamp 0
transform 1 0 16836 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_195
timestamp 0
transform 1 0 19596 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_196
timestamp 0
transform 1 0 22356 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_197
timestamp 0
transform 1 0 25116 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp 0
transform 1 0 27876 0 -1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_199
timestamp 0
transform 1 0 4416 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_200
timestamp 0
transform 1 0 7176 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_201
timestamp 0
transform 1 0 9936 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_202
timestamp 0
transform 1 0 12696 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp 0
transform 1 0 15456 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_204
timestamp 0
transform 1 0 18216 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_205
timestamp 0
transform 1 0 20976 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_206
timestamp 0
transform 1 0 23736 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_207
timestamp 0
transform 1 0 26496 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_208
timestamp 0
transform 1 0 29256 0 1 8704
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_209
timestamp 0
transform 1 0 5796 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_210
timestamp 0
transform 1 0 8556 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_211
timestamp 0
transform 1 0 11316 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_212
timestamp 0
transform 1 0 14076 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_213
timestamp 0
transform 1 0 16836 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_214
timestamp 0
transform 1 0 19596 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_215
timestamp 0
transform 1 0 22356 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_216
timestamp 0
transform 1 0 25116 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_217
timestamp 0
transform 1 0 27876 0 -1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_218
timestamp 0
transform 1 0 4416 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_219
timestamp 0
transform 1 0 7176 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_220
timestamp 0
transform 1 0 9936 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_221
timestamp 0
transform 1 0 12696 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_222
timestamp 0
transform 1 0 15456 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_223
timestamp 0
transform 1 0 18216 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_224
timestamp 0
transform 1 0 20976 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_225
timestamp 0
transform 1 0 23736 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_226
timestamp 0
transform 1 0 26496 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_227
timestamp 0
transform 1 0 29256 0 1 9248
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_228
timestamp 0
transform 1 0 5796 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_229
timestamp 0
transform 1 0 8556 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_230
timestamp 0
transform 1 0 11316 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_231
timestamp 0
transform 1 0 14076 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_232
timestamp 0
transform 1 0 16836 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_233
timestamp 0
transform 1 0 19596 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_234
timestamp 0
transform 1 0 22356 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_235
timestamp 0
transform 1 0 25116 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_236
timestamp 0
transform 1 0 27876 0 -1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_237
timestamp 0
transform 1 0 4416 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_238
timestamp 0
transform 1 0 7176 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_239
timestamp 0
transform 1 0 9936 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_240
timestamp 0
transform 1 0 12696 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_241
timestamp 0
transform 1 0 15456 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_242
timestamp 0
transform 1 0 18216 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_243
timestamp 0
transform 1 0 20976 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_244
timestamp 0
transform 1 0 23736 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_245
timestamp 0
transform 1 0 26496 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_246
timestamp 0
transform 1 0 29256 0 1 9792
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_247
timestamp 0
transform 1 0 5796 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_248
timestamp 0
transform 1 0 8556 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_249
timestamp 0
transform 1 0 11316 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_250
timestamp 0
transform 1 0 14076 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_251
timestamp 0
transform 1 0 16836 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_252
timestamp 0
transform 1 0 19596 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_253
timestamp 0
transform 1 0 22356 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_254
timestamp 0
transform 1 0 25116 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_255
timestamp 0
transform 1 0 27876 0 -1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_256
timestamp 0
transform 1 0 4416 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_257
timestamp 0
transform 1 0 7176 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_258
timestamp 0
transform 1 0 9936 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_259
timestamp 0
transform 1 0 12696 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_260
timestamp 0
transform 1 0 15456 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_261
timestamp 0
transform 1 0 18216 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_262
timestamp 0
transform 1 0 20976 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_263
timestamp 0
transform 1 0 23736 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_264
timestamp 0
transform 1 0 26496 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_265
timestamp 0
transform 1 0 29256 0 1 10336
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_266
timestamp 0
transform 1 0 5796 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_267
timestamp 0
transform 1 0 8556 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_268
timestamp 0
transform 1 0 11316 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_269
timestamp 0
transform 1 0 14076 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_270
timestamp 0
transform 1 0 16836 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_271
timestamp 0
transform 1 0 19596 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_272
timestamp 0
transform 1 0 22356 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_273
timestamp 0
transform 1 0 25116 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_274
timestamp 0
transform 1 0 27876 0 -1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_275
timestamp 0
transform 1 0 4416 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_276
timestamp 0
transform 1 0 7176 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_277
timestamp 0
transform 1 0 9936 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_278
timestamp 0
transform 1 0 12696 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_279
timestamp 0
transform 1 0 15456 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_280
timestamp 0
transform 1 0 18216 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_281
timestamp 0
transform 1 0 20976 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_282
timestamp 0
transform 1 0 23736 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_283
timestamp 0
transform 1 0 26496 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_284
timestamp 0
transform 1 0 29256 0 1 10880
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_285
timestamp 0
transform 1 0 5796 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_286
timestamp 0
transform 1 0 8556 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_287
timestamp 0
transform 1 0 11316 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_288
timestamp 0
transform 1 0 14076 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_289
timestamp 0
transform 1 0 16836 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_290
timestamp 0
transform 1 0 19596 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_291
timestamp 0
transform 1 0 22356 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_292
timestamp 0
transform 1 0 25116 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_293
timestamp 0
transform 1 0 27876 0 -1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_294
timestamp 0
transform 1 0 4416 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_295
timestamp 0
transform 1 0 7176 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_296
timestamp 0
transform 1 0 9936 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_297
timestamp 0
transform 1 0 12696 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_298
timestamp 0
transform 1 0 15456 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_299
timestamp 0
transform 1 0 18216 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_300
timestamp 0
transform 1 0 20976 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_301
timestamp 0
transform 1 0 23736 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_302
timestamp 0
transform 1 0 26496 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_303
timestamp 0
transform 1 0 29256 0 1 11424
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_304
timestamp 0
transform 1 0 5796 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_305
timestamp 0
transform 1 0 8556 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_306
timestamp 0
transform 1 0 11316 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_307
timestamp 0
transform 1 0 14076 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_308
timestamp 0
transform 1 0 16836 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_309
timestamp 0
transform 1 0 19596 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_310
timestamp 0
transform 1 0 22356 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_311
timestamp 0
transform 1 0 25116 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_312
timestamp 0
transform 1 0 27876 0 -1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_313
timestamp 0
transform 1 0 4416 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_314
timestamp 0
transform 1 0 7176 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_315
timestamp 0
transform 1 0 9936 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_316
timestamp 0
transform 1 0 12696 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_317
timestamp 0
transform 1 0 15456 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_318
timestamp 0
transform 1 0 18216 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_319
timestamp 0
transform 1 0 20976 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_320
timestamp 0
transform 1 0 23736 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_321
timestamp 0
transform 1 0 26496 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_322
timestamp 0
transform 1 0 29256 0 1 11968
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_323
timestamp 0
transform 1 0 5796 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_324
timestamp 0
transform 1 0 8556 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_325
timestamp 0
transform 1 0 11316 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_326
timestamp 0
transform 1 0 14076 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_327
timestamp 0
transform 1 0 16836 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_328
timestamp 0
transform 1 0 19596 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_329
timestamp 0
transform 1 0 22356 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_330
timestamp 0
transform 1 0 25116 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_331
timestamp 0
transform 1 0 27876 0 -1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_332
timestamp 0
transform 1 0 4416 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_333
timestamp 0
transform 1 0 7176 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_334
timestamp 0
transform 1 0 9936 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_335
timestamp 0
transform 1 0 12696 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_336
timestamp 0
transform 1 0 15456 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_337
timestamp 0
transform 1 0 18216 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_338
timestamp 0
transform 1 0 20976 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_339
timestamp 0
transform 1 0 23736 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_340
timestamp 0
transform 1 0 26496 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_341
timestamp 0
transform 1 0 29256 0 1 12512
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_342
timestamp 0
transform 1 0 5796 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_343
timestamp 0
transform 1 0 8556 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_344
timestamp 0
transform 1 0 11316 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_345
timestamp 0
transform 1 0 14076 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_346
timestamp 0
transform 1 0 16836 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_347
timestamp 0
transform 1 0 19596 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_348
timestamp 0
transform 1 0 22356 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_349
timestamp 0
transform 1 0 25116 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_350
timestamp 0
transform 1 0 27876 0 -1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_351
timestamp 0
transform 1 0 4416 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_352
timestamp 0
transform 1 0 7176 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_353
timestamp 0
transform 1 0 9936 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_354
timestamp 0
transform 1 0 12696 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_355
timestamp 0
transform 1 0 15456 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_356
timestamp 0
transform 1 0 18216 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_357
timestamp 0
transform 1 0 20976 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_358
timestamp 0
transform 1 0 23736 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_359
timestamp 0
transform 1 0 26496 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_360
timestamp 0
transform 1 0 29256 0 1 13056
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_361
timestamp 0
transform 1 0 5796 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_362
timestamp 0
transform 1 0 8556 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_363
timestamp 0
transform 1 0 11316 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_364
timestamp 0
transform 1 0 14076 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_365
timestamp 0
transform 1 0 16836 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_366
timestamp 0
transform 1 0 19596 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_367
timestamp 0
transform 1 0 22356 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_368
timestamp 0
transform 1 0 25116 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_369
timestamp 0
transform 1 0 27876 0 -1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_370
timestamp 0
transform 1 0 4416 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_371
timestamp 0
transform 1 0 7176 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_372
timestamp 0
transform 1 0 9936 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_373
timestamp 0
transform 1 0 12696 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_374
timestamp 0
transform 1 0 15456 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_375
timestamp 0
transform 1 0 18216 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_376
timestamp 0
transform 1 0 20976 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_377
timestamp 0
transform 1 0 23736 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_378
timestamp 0
transform 1 0 26496 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_379
timestamp 0
transform 1 0 29256 0 1 13600
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_380
timestamp 0
transform 1 0 5796 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_381
timestamp 0
transform 1 0 8556 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_382
timestamp 0
transform 1 0 11316 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_383
timestamp 0
transform 1 0 14076 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_384
timestamp 0
transform 1 0 16836 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_385
timestamp 0
transform 1 0 19596 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_386
timestamp 0
transform 1 0 22356 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_387
timestamp 0
transform 1 0 25116 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_388
timestamp 0
transform 1 0 27876 0 -1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_389
timestamp 0
transform 1 0 4416 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_390
timestamp 0
transform 1 0 7176 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_391
timestamp 0
transform 1 0 9936 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_392
timestamp 0
transform 1 0 12696 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_393
timestamp 0
transform 1 0 15456 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_394
timestamp 0
transform 1 0 18216 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_395
timestamp 0
transform 1 0 20976 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_396
timestamp 0
transform 1 0 23736 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_397
timestamp 0
transform 1 0 26496 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_398
timestamp 0
transform 1 0 29256 0 1 14144
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_399
timestamp 0
transform 1 0 5796 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_400
timestamp 0
transform 1 0 8556 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_401
timestamp 0
transform 1 0 11316 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_402
timestamp 0
transform 1 0 14076 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_403
timestamp 0
transform 1 0 16836 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_404
timestamp 0
transform 1 0 19596 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_405
timestamp 0
transform 1 0 22356 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_406
timestamp 0
transform 1 0 25116 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_407
timestamp 0
transform 1 0 27876 0 -1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_408
timestamp 0
transform 1 0 4416 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_409
timestamp 0
transform 1 0 7176 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_410
timestamp 0
transform 1 0 9936 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_411
timestamp 0
transform 1 0 12696 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_412
timestamp 0
transform 1 0 15456 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_413
timestamp 0
transform 1 0 18216 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_414
timestamp 0
transform 1 0 20976 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_415
timestamp 0
transform 1 0 23736 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_416
timestamp 0
transform 1 0 26496 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_417
timestamp 0
transform 1 0 29256 0 1 14688
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_418
timestamp 0
transform 1 0 5796 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_419
timestamp 0
transform 1 0 8556 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_420
timestamp 0
transform 1 0 11316 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_421
timestamp 0
transform 1 0 14076 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_422
timestamp 0
transform 1 0 16836 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_423
timestamp 0
transform 1 0 19596 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_424
timestamp 0
transform 1 0 22356 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_425
timestamp 0
transform 1 0 25116 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_426
timestamp 0
transform 1 0 27876 0 -1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_427
timestamp 0
transform 1 0 4416 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_428
timestamp 0
transform 1 0 7176 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_429
timestamp 0
transform 1 0 9936 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_430
timestamp 0
transform 1 0 12696 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_431
timestamp 0
transform 1 0 15456 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_432
timestamp 0
transform 1 0 18216 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_433
timestamp 0
transform 1 0 20976 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_434
timestamp 0
transform 1 0 23736 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_435
timestamp 0
transform 1 0 26496 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_436
timestamp 0
transform 1 0 29256 0 1 15232
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_437
timestamp 0
transform 1 0 5796 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_438
timestamp 0
transform 1 0 8556 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_439
timestamp 0
transform 1 0 11316 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_440
timestamp 0
transform 1 0 14076 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_441
timestamp 0
transform 1 0 16836 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_442
timestamp 0
transform 1 0 19596 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_443
timestamp 0
transform 1 0 22356 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_444
timestamp 0
transform 1 0 25116 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_445
timestamp 0
transform 1 0 27876 0 -1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_446
timestamp 0
transform 1 0 4416 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_447
timestamp 0
transform 1 0 7176 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_448
timestamp 0
transform 1 0 9936 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_449
timestamp 0
transform 1 0 12696 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_450
timestamp 0
transform 1 0 15456 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_451
timestamp 0
transform 1 0 18216 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_452
timestamp 0
transform 1 0 20976 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_453
timestamp 0
transform 1 0 23736 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_454
timestamp 0
transform 1 0 26496 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_455
timestamp 0
transform 1 0 29256 0 1 15776
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_456
timestamp 0
transform 1 0 5796 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_457
timestamp 0
transform 1 0 8556 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_458
timestamp 0
transform 1 0 11316 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_459
timestamp 0
transform 1 0 14076 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_460
timestamp 0
transform 1 0 16836 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_461
timestamp 0
transform 1 0 19596 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_462
timestamp 0
transform 1 0 22356 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_463
timestamp 0
transform 1 0 25116 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_464
timestamp 0
transform 1 0 27876 0 -1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_465
timestamp 0
transform 1 0 4416 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_466
timestamp 0
transform 1 0 7176 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_467
timestamp 0
transform 1 0 9936 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_468
timestamp 0
transform 1 0 12696 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_469
timestamp 0
transform 1 0 15456 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_470
timestamp 0
transform 1 0 18216 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_471
timestamp 0
transform 1 0 20976 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_472
timestamp 0
transform 1 0 23736 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_473
timestamp 0
transform 1 0 26496 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_474
timestamp 0
transform 1 0 29256 0 1 16320
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_475
timestamp 0
transform 1 0 5796 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_476
timestamp 0
transform 1 0 8556 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_477
timestamp 0
transform 1 0 11316 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_478
timestamp 0
transform 1 0 14076 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_479
timestamp 0
transform 1 0 16836 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_480
timestamp 0
transform 1 0 19596 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_481
timestamp 0
transform 1 0 22356 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_482
timestamp 0
transform 1 0 25116 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_483
timestamp 0
transform 1 0 27876 0 -1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_484
timestamp 0
transform 1 0 4416 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_485
timestamp 0
transform 1 0 7176 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_486
timestamp 0
transform 1 0 9936 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_487
timestamp 0
transform 1 0 12696 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_488
timestamp 0
transform 1 0 15456 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_489
timestamp 0
transform 1 0 18216 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_490
timestamp 0
transform 1 0 20976 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_491
timestamp 0
transform 1 0 23736 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_492
timestamp 0
transform 1 0 26496 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_493
timestamp 0
transform 1 0 29256 0 1 16864
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_494
timestamp 0
transform 1 0 5796 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_495
timestamp 0
transform 1 0 8556 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_496
timestamp 0
transform 1 0 11316 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_497
timestamp 0
transform 1 0 14076 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_498
timestamp 0
transform 1 0 16836 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_499
timestamp 0
transform 1 0 19596 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_500
timestamp 0
transform 1 0 22356 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_501
timestamp 0
transform 1 0 25116 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_502
timestamp 0
transform 1 0 27876 0 -1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_503
timestamp 0
transform 1 0 4416 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_504
timestamp 0
transform 1 0 7176 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_505
timestamp 0
transform 1 0 9936 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_506
timestamp 0
transform 1 0 12696 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_507
timestamp 0
transform 1 0 15456 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_508
timestamp 0
transform 1 0 18216 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_509
timestamp 0
transform 1 0 20976 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_510
timestamp 0
transform 1 0 23736 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_511
timestamp 0
transform 1 0 26496 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_512
timestamp 0
transform 1 0 29256 0 1 17408
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_513
timestamp 0
transform 1 0 5796 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_514
timestamp 0
transform 1 0 8556 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_515
timestamp 0
transform 1 0 11316 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_516
timestamp 0
transform 1 0 14076 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_517
timestamp 0
transform 1 0 16836 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_518
timestamp 0
transform 1 0 19596 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_519
timestamp 0
transform 1 0 22356 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_520
timestamp 0
transform 1 0 25116 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_521
timestamp 0
transform 1 0 27876 0 -1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_522
timestamp 0
transform 1 0 4416 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_523
timestamp 0
transform 1 0 7176 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_524
timestamp 0
transform 1 0 9936 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_525
timestamp 0
transform 1 0 12696 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_526
timestamp 0
transform 1 0 15456 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_527
timestamp 0
transform 1 0 18216 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_528
timestamp 0
transform 1 0 20976 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_529
timestamp 0
transform 1 0 23736 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_530
timestamp 0
transform 1 0 26496 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_531
timestamp 0
transform 1 0 29256 0 1 17952
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_532
timestamp 0
transform 1 0 5796 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_533
timestamp 0
transform 1 0 8556 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_534
timestamp 0
transform 1 0 11316 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_535
timestamp 0
transform 1 0 14076 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_536
timestamp 0
transform 1 0 16836 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_537
timestamp 0
transform 1 0 19596 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_538
timestamp 0
transform 1 0 22356 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_539
timestamp 0
transform 1 0 25116 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_540
timestamp 0
transform 1 0 27876 0 -1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_541
timestamp 0
transform 1 0 4416 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_542
timestamp 0
transform 1 0 7176 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_543
timestamp 0
transform 1 0 9936 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_544
timestamp 0
transform 1 0 12696 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_545
timestamp 0
transform 1 0 15456 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_546
timestamp 0
transform 1 0 18216 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_547
timestamp 0
transform 1 0 20976 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_548
timestamp 0
transform 1 0 23736 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_549
timestamp 0
transform 1 0 26496 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_550
timestamp 0
transform 1 0 29256 0 1 18496
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_551
timestamp 0
transform 1 0 5796 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_552
timestamp 0
transform 1 0 8556 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_553
timestamp 0
transform 1 0 11316 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_554
timestamp 0
transform 1 0 14076 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_555
timestamp 0
transform 1 0 16836 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_556
timestamp 0
transform 1 0 19596 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_557
timestamp 0
transform 1 0 22356 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_558
timestamp 0
transform 1 0 25116 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_559
timestamp 0
transform 1 0 27876 0 -1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_560
timestamp 0
transform 1 0 4416 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_561
timestamp 0
transform 1 0 7176 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_562
timestamp 0
transform 1 0 9936 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_563
timestamp 0
transform 1 0 12696 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_564
timestamp 0
transform 1 0 15456 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_565
timestamp 0
transform 1 0 18216 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_566
timestamp 0
transform 1 0 20976 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_567
timestamp 0
transform 1 0 23736 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_568
timestamp 0
transform 1 0 26496 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_569
timestamp 0
transform 1 0 29256 0 1 19040
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_570
timestamp 0
transform 1 0 5796 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_571
timestamp 0
transform 1 0 8556 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_572
timestamp 0
transform 1 0 11316 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_573
timestamp 0
transform 1 0 14076 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_574
timestamp 0
transform 1 0 16836 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_575
timestamp 0
transform 1 0 19596 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_576
timestamp 0
transform 1 0 22356 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_577
timestamp 0
transform 1 0 25116 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_578
timestamp 0
transform 1 0 27876 0 -1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_579
timestamp 0
transform 1 0 4416 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_580
timestamp 0
transform 1 0 7176 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_581
timestamp 0
transform 1 0 9936 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_582
timestamp 0
transform 1 0 12696 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_583
timestamp 0
transform 1 0 15456 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_584
timestamp 0
transform 1 0 18216 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_585
timestamp 0
transform 1 0 20976 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_586
timestamp 0
transform 1 0 23736 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_587
timestamp 0
transform 1 0 26496 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_588
timestamp 0
transform 1 0 29256 0 1 19584
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_589
timestamp 0
transform 1 0 5796 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_590
timestamp 0
transform 1 0 8556 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_591
timestamp 0
transform 1 0 11316 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_592
timestamp 0
transform 1 0 14076 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_593
timestamp 0
transform 1 0 16836 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_594
timestamp 0
transform 1 0 19596 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_595
timestamp 0
transform 1 0 22356 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_596
timestamp 0
transform 1 0 25116 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_597
timestamp 0
transform 1 0 27876 0 -1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_598
timestamp 0
transform 1 0 4416 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_599
timestamp 0
transform 1 0 7176 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_600
timestamp 0
transform 1 0 9936 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_601
timestamp 0
transform 1 0 12696 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_602
timestamp 0
transform 1 0 15456 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_603
timestamp 0
transform 1 0 18216 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_604
timestamp 0
transform 1 0 20976 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_605
timestamp 0
transform 1 0 23736 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_606
timestamp 0
transform 1 0 26496 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_607
timestamp 0
transform 1 0 29256 0 1 20128
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_608
timestamp 0
transform 1 0 5796 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_609
timestamp 0
transform 1 0 8556 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_610
timestamp 0
transform 1 0 11316 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_611
timestamp 0
transform 1 0 14076 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_612
timestamp 0
transform 1 0 16836 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_613
timestamp 0
transform 1 0 19596 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_614
timestamp 0
transform 1 0 22356 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_615
timestamp 0
transform 1 0 25116 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_616
timestamp 0
transform 1 0 27876 0 -1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_617
timestamp 0
transform 1 0 4416 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_618
timestamp 0
transform 1 0 7176 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_619
timestamp 0
transform 1 0 9936 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_620
timestamp 0
transform 1 0 12696 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_621
timestamp 0
transform 1 0 15456 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_622
timestamp 0
transform 1 0 18216 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_623
timestamp 0
transform 1 0 20976 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_624
timestamp 0
transform 1 0 23736 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_625
timestamp 0
transform 1 0 26496 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_626
timestamp 0
transform 1 0 29256 0 1 20672
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_627
timestamp 0
transform 1 0 5796 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_628
timestamp 0
transform 1 0 8556 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_629
timestamp 0
transform 1 0 11316 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_630
timestamp 0
transform 1 0 14076 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_631
timestamp 0
transform 1 0 16836 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_632
timestamp 0
transform 1 0 19596 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_633
timestamp 0
transform 1 0 22356 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_634
timestamp 0
transform 1 0 25116 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_635
timestamp 0
transform 1 0 27876 0 -1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_636
timestamp 0
transform 1 0 4416 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_637
timestamp 0
transform 1 0 7176 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_638
timestamp 0
transform 1 0 9936 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_639
timestamp 0
transform 1 0 12696 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_640
timestamp 0
transform 1 0 15456 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_641
timestamp 0
transform 1 0 18216 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_642
timestamp 0
transform 1 0 20976 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_643
timestamp 0
transform 1 0 23736 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_644
timestamp 0
transform 1 0 26496 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_645
timestamp 0
transform 1 0 29256 0 1 21216
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_646
timestamp 0
transform 1 0 5796 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_647
timestamp 0
transform 1 0 8556 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_648
timestamp 0
transform 1 0 11316 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_649
timestamp 0
transform 1 0 14076 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_650
timestamp 0
transform 1 0 16836 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_651
timestamp 0
transform 1 0 19596 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_652
timestamp 0
transform 1 0 22356 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_653
timestamp 0
transform 1 0 25116 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_654
timestamp 0
transform 1 0 27876 0 -1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_655
timestamp 0
transform 1 0 4416 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_656
timestamp 0
transform 1 0 7176 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_657
timestamp 0
transform 1 0 9936 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_658
timestamp 0
transform 1 0 12696 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_659
timestamp 0
transform 1 0 15456 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_660
timestamp 0
transform 1 0 18216 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_661
timestamp 0
transform 1 0 20976 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_662
timestamp 0
transform 1 0 23736 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_663
timestamp 0
transform 1 0 26496 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_664
timestamp 0
transform 1 0 29256 0 1 21760
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_665
timestamp 0
transform 1 0 5796 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_666
timestamp 0
transform 1 0 8556 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_667
timestamp 0
transform 1 0 11316 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_668
timestamp 0
transform 1 0 14076 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_669
timestamp 0
transform 1 0 16836 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_670
timestamp 0
transform 1 0 19596 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_671
timestamp 0
transform 1 0 22356 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_672
timestamp 0
transform 1 0 25116 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_673
timestamp 0
transform 1 0 27876 0 -1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_674
timestamp 0
transform 1 0 4416 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_675
timestamp 0
transform 1 0 7176 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_676
timestamp 0
transform 1 0 9936 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_677
timestamp 0
transform 1 0 12696 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_678
timestamp 0
transform 1 0 15456 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_679
timestamp 0
transform 1 0 18216 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_680
timestamp 0
transform 1 0 20976 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_681
timestamp 0
transform 1 0 23736 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_682
timestamp 0
transform 1 0 26496 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_683
timestamp 0
transform 1 0 29256 0 1 22304
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_684
timestamp 0
transform 1 0 5796 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_685
timestamp 0
transform 1 0 8556 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_686
timestamp 0
transform 1 0 11316 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_687
timestamp 0
transform 1 0 14076 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_688
timestamp 0
transform 1 0 16836 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_689
timestamp 0
transform 1 0 19596 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_690
timestamp 0
transform 1 0 22356 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_691
timestamp 0
transform 1 0 25116 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_692
timestamp 0
transform 1 0 27876 0 -1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_693
timestamp 0
transform 1 0 4416 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_694
timestamp 0
transform 1 0 7176 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_695
timestamp 0
transform 1 0 9936 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_696
timestamp 0
transform 1 0 12696 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_697
timestamp 0
transform 1 0 15456 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_698
timestamp 0
transform 1 0 18216 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_699
timestamp 0
transform 1 0 20976 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_700
timestamp 0
transform 1 0 23736 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_701
timestamp 0
transform 1 0 26496 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_702
timestamp 0
transform 1 0 29256 0 1 22848
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_703
timestamp 0
transform 1 0 5796 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_704
timestamp 0
transform 1 0 8556 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_705
timestamp 0
transform 1 0 11316 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_706
timestamp 0
transform 1 0 14076 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_707
timestamp 0
transform 1 0 16836 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_708
timestamp 0
transform 1 0 19596 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_709
timestamp 0
transform 1 0 22356 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_710
timestamp 0
transform 1 0 25116 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_711
timestamp 0
transform 1 0 27876 0 -1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_712
timestamp 0
transform 1 0 4416 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_713
timestamp 0
transform 1 0 7176 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_714
timestamp 0
transform 1 0 9936 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_715
timestamp 0
transform 1 0 12696 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_716
timestamp 0
transform 1 0 15456 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_717
timestamp 0
transform 1 0 18216 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_718
timestamp 0
transform 1 0 20976 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_719
timestamp 0
transform 1 0 23736 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_720
timestamp 0
transform 1 0 26496 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_721
timestamp 0
transform 1 0 29256 0 1 23392
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_722
timestamp 0
transform 1 0 5796 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_723
timestamp 0
transform 1 0 8556 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_724
timestamp 0
transform 1 0 11316 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_725
timestamp 0
transform 1 0 14076 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_726
timestamp 0
transform 1 0 16836 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_727
timestamp 0
transform 1 0 19596 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_728
timestamp 0
transform 1 0 22356 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_729
timestamp 0
transform 1 0 25116 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_730
timestamp 0
transform 1 0 27876 0 -1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_731
timestamp 0
transform 1 0 4416 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_732
timestamp 0
transform 1 0 7176 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_733
timestamp 0
transform 1 0 9936 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_734
timestamp 0
transform 1 0 12696 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_735
timestamp 0
transform 1 0 15456 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_736
timestamp 0
transform 1 0 18216 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_737
timestamp 0
transform 1 0 20976 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_738
timestamp 0
transform 1 0 23736 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_739
timestamp 0
transform 1 0 26496 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_740
timestamp 0
transform 1 0 29256 0 1 23936
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_741
timestamp 0
transform 1 0 5796 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_742
timestamp 0
transform 1 0 8556 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_743
timestamp 0
transform 1 0 11316 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_744
timestamp 0
transform 1 0 14076 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_745
timestamp 0
transform 1 0 16836 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_746
timestamp 0
transform 1 0 19596 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_747
timestamp 0
transform 1 0 22356 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_748
timestamp 0
transform 1 0 25116 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_749
timestamp 0
transform 1 0 27876 0 -1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_750
timestamp 0
transform 1 0 4416 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_751
timestamp 0
transform 1 0 7176 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_752
timestamp 0
transform 1 0 9936 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_753
timestamp 0
transform 1 0 12696 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_754
timestamp 0
transform 1 0 15456 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_755
timestamp 0
transform 1 0 18216 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_756
timestamp 0
transform 1 0 20976 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_757
timestamp 0
transform 1 0 23736 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_758
timestamp 0
transform 1 0 26496 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_759
timestamp 0
transform 1 0 29256 0 1 24480
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_760
timestamp 0
transform 1 0 5796 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_761
timestamp 0
transform 1 0 8556 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_762
timestamp 0
transform 1 0 11316 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_763
timestamp 0
transform 1 0 14076 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_764
timestamp 0
transform 1 0 16836 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_765
timestamp 0
transform 1 0 19596 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_766
timestamp 0
transform 1 0 22356 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_767
timestamp 0
transform 1 0 25116 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_768
timestamp 0
transform 1 0 27876 0 -1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_769
timestamp 0
transform 1 0 4416 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_770
timestamp 0
transform 1 0 7176 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_771
timestamp 0
transform 1 0 9936 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_772
timestamp 0
transform 1 0 12696 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_773
timestamp 0
transform 1 0 15456 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_774
timestamp 0
transform 1 0 18216 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_775
timestamp 0
transform 1 0 20976 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_776
timestamp 0
transform 1 0 23736 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_777
timestamp 0
transform 1 0 26496 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_778
timestamp 0
transform 1 0 29256 0 1 25024
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_779
timestamp 0
transform 1 0 5796 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_780
timestamp 0
transform 1 0 8556 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_781
timestamp 0
transform 1 0 11316 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_782
timestamp 0
transform 1 0 14076 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_783
timestamp 0
transform 1 0 16836 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_784
timestamp 0
transform 1 0 19596 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_785
timestamp 0
transform 1 0 22356 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_786
timestamp 0
transform 1 0 25116 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_787
timestamp 0
transform 1 0 27876 0 -1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_788
timestamp 0
transform 1 0 4416 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_789
timestamp 0
transform 1 0 7176 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_790
timestamp 0
transform 1 0 9936 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_791
timestamp 0
transform 1 0 12696 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_792
timestamp 0
transform 1 0 15456 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_793
timestamp 0
transform 1 0 18216 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_794
timestamp 0
transform 1 0 20976 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_795
timestamp 0
transform 1 0 23736 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_796
timestamp 0
transform 1 0 26496 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_797
timestamp 0
transform 1 0 29256 0 1 25568
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_798
timestamp 0
transform 1 0 5796 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_799
timestamp 0
transform 1 0 8556 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_800
timestamp 0
transform 1 0 11316 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_801
timestamp 0
transform 1 0 14076 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_802
timestamp 0
transform 1 0 16836 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_803
timestamp 0
transform 1 0 19596 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_804
timestamp 0
transform 1 0 22356 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_805
timestamp 0
transform 1 0 25116 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_806
timestamp 0
transform 1 0 27876 0 -1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_807
timestamp 0
transform 1 0 4416 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_808
timestamp 0
transform 1 0 7176 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_809
timestamp 0
transform 1 0 9936 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_810
timestamp 0
transform 1 0 12696 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_811
timestamp 0
transform 1 0 15456 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_812
timestamp 0
transform 1 0 18216 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_813
timestamp 0
transform 1 0 20976 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_814
timestamp 0
transform 1 0 23736 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_815
timestamp 0
transform 1 0 26496 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_816
timestamp 0
transform 1 0 29256 0 1 26112
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_817
timestamp 0
transform 1 0 5796 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_818
timestamp 0
transform 1 0 8556 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_819
timestamp 0
transform 1 0 11316 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_820
timestamp 0
transform 1 0 14076 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_821
timestamp 0
transform 1 0 16836 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_822
timestamp 0
transform 1 0 19596 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_823
timestamp 0
transform 1 0 22356 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_824
timestamp 0
transform 1 0 25116 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_825
timestamp 0
transform 1 0 27876 0 -1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_826
timestamp 0
transform 1 0 4416 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_827
timestamp 0
transform 1 0 7176 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_828
timestamp 0
transform 1 0 9936 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_829
timestamp 0
transform 1 0 12696 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_830
timestamp 0
transform 1 0 15456 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_831
timestamp 0
transform 1 0 18216 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_832
timestamp 0
transform 1 0 20976 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_833
timestamp 0
transform 1 0 23736 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_834
timestamp 0
transform 1 0 26496 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_835
timestamp 0
transform 1 0 29256 0 1 26656
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_836
timestamp 0
transform 1 0 5796 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_837
timestamp 0
transform 1 0 8556 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_838
timestamp 0
transform 1 0 11316 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_839
timestamp 0
transform 1 0 14076 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_840
timestamp 0
transform 1 0 16836 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_841
timestamp 0
transform 1 0 19596 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_842
timestamp 0
transform 1 0 22356 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_843
timestamp 0
transform 1 0 25116 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_844
timestamp 0
transform 1 0 27876 0 -1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_845
timestamp 0
transform 1 0 4416 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_846
timestamp 0
transform 1 0 7176 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_847
timestamp 0
transform 1 0 9936 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_848
timestamp 0
transform 1 0 12696 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_849
timestamp 0
transform 1 0 15456 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_850
timestamp 0
transform 1 0 18216 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_851
timestamp 0
transform 1 0 20976 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_852
timestamp 0
transform 1 0 23736 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_853
timestamp 0
transform 1 0 26496 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_854
timestamp 0
transform 1 0 29256 0 1 27200
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_855
timestamp 0
transform 1 0 5796 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_856
timestamp 0
transform 1 0 8556 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_857
timestamp 0
transform 1 0 11316 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_858
timestamp 0
transform 1 0 14076 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_859
timestamp 0
transform 1 0 16836 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_860
timestamp 0
transform 1 0 19596 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_861
timestamp 0
transform 1 0 22356 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_862
timestamp 0
transform 1 0 25116 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_863
timestamp 0
transform 1 0 27876 0 -1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_864
timestamp 0
transform 1 0 4416 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_865
timestamp 0
transform 1 0 7176 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_866
timestamp 0
transform 1 0 9936 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_867
timestamp 0
transform 1 0 12696 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_868
timestamp 0
transform 1 0 15456 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_869
timestamp 0
transform 1 0 18216 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_870
timestamp 0
transform 1 0 20976 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_871
timestamp 0
transform 1 0 23736 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_872
timestamp 0
transform 1 0 26496 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_873
timestamp 0
transform 1 0 29256 0 1 27744
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_874
timestamp 0
transform 1 0 5796 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_875
timestamp 0
transform 1 0 8556 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_876
timestamp 0
transform 1 0 11316 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_877
timestamp 0
transform 1 0 14076 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_878
timestamp 0
transform 1 0 16836 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_879
timestamp 0
transform 1 0 19596 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_880
timestamp 0
transform 1 0 22356 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_881
timestamp 0
transform 1 0 25116 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_882
timestamp 0
transform 1 0 27876 0 -1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_883
timestamp 0
transform 1 0 4416 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_884
timestamp 0
transform 1 0 7176 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_885
timestamp 0
transform 1 0 9936 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_886
timestamp 0
transform 1 0 12696 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_887
timestamp 0
transform 1 0 15456 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_888
timestamp 0
transform 1 0 18216 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_889
timestamp 0
transform 1 0 20976 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_890
timestamp 0
transform 1 0 23736 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_891
timestamp 0
transform 1 0 26496 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_892
timestamp 0
transform 1 0 29256 0 1 28288
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_893
timestamp 0
transform 1 0 5796 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_894
timestamp 0
transform 1 0 8556 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_895
timestamp 0
transform 1 0 11316 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_896
timestamp 0
transform 1 0 14076 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_897
timestamp 0
transform 1 0 16836 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_898
timestamp 0
transform 1 0 19596 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_899
timestamp 0
transform 1 0 22356 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_900
timestamp 0
transform 1 0 25116 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_901
timestamp 0
transform 1 0 27876 0 -1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_902
timestamp 0
transform 1 0 4416 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_903
timestamp 0
transform 1 0 7176 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_904
timestamp 0
transform 1 0 9936 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_905
timestamp 0
transform 1 0 12696 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_906
timestamp 0
transform 1 0 15456 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_907
timestamp 0
transform 1 0 18216 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_908
timestamp 0
transform 1 0 20976 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_909
timestamp 0
transform 1 0 23736 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_910
timestamp 0
transform 1 0 26496 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_911
timestamp 0
transform 1 0 29256 0 1 28832
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_912
timestamp 0
transform 1 0 5796 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_913
timestamp 0
transform 1 0 8556 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_914
timestamp 0
transform 1 0 11316 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_915
timestamp 0
transform 1 0 14076 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_916
timestamp 0
transform 1 0 16836 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_917
timestamp 0
transform 1 0 19596 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_918
timestamp 0
transform 1 0 22356 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_919
timestamp 0
transform 1 0 25116 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_920
timestamp 0
transform 1 0 27876 0 -1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_921
timestamp 0
transform 1 0 4416 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_922
timestamp 0
transform 1 0 7176 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_923
timestamp 0
transform 1 0 9936 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_924
timestamp 0
transform 1 0 12696 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_925
timestamp 0
transform 1 0 15456 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_926
timestamp 0
transform 1 0 18216 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_927
timestamp 0
transform 1 0 20976 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_928
timestamp 0
transform 1 0 23736 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_929
timestamp 0
transform 1 0 26496 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_930
timestamp 0
transform 1 0 29256 0 1 29376
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_931
timestamp 0
transform 1 0 4416 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_932
timestamp 0
transform 1 0 5796 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_933
timestamp 0
transform 1 0 7176 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_934
timestamp 0
transform 1 0 8556 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_935
timestamp 0
transform 1 0 9936 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_936
timestamp 0
transform 1 0 11316 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_937
timestamp 0
transform 1 0 12696 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_938
timestamp 0
transform 1 0 14076 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_939
timestamp 0
transform 1 0 15456 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_940
timestamp 0
transform 1 0 16836 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_941
timestamp 0
transform 1 0 18216 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_942
timestamp 0
transform 1 0 19596 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_943
timestamp 0
transform 1 0 20976 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_944
timestamp 0
transform 1 0 22356 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_945
timestamp 0
transform 1 0 23736 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_946
timestamp 0
transform 1 0 25116 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_947
timestamp 0
transform 1 0 26496 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_948
timestamp 0
transform 1 0 27876 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_949
timestamp 0
transform 1 0 29256 0 -1 29920
box 0 -24 46 296
use sky130_fd_sc_hd__clkbuf_4  wire1
timestamp 0
transform 1 0 16284 0 1 23936
box 0 -24 276 296
<< labels >>
flabel metal3 s 32920 15251 33000 15281 0 FreeSans 240 0 0 0 BE
port 0 nsew signal output
flabel metal2 s 15748 0 15762 48 0 FreeSans 112 90 0 0 FE
port 1 nsew signal output
flabel metal2 s 11884 0 11898 48 0 FreeSans 112 90 0 0 OE
port 2 nsew signal output
flabel metal2 s 5536 0 5550 48 0 FreeSans 112 90 0 0 SysClk
port 3 nsew signal input
flabel metal2 s 7836 0 7850 48 0 FreeSans 112 90 0 0 baud_selector[0]
port 4 nsew signal input
flabel metal2 s 7744 0 7758 48 0 FreeSans 112 90 0 0 baud_selector[1]
port 5 nsew signal input
flabel metal2 s 18784 0 18798 48 0 FreeSans 112 90 0 0 data_in[0]
port 6 nsew signal input
flabel metal2 s 22832 32952 22846 33000 0 FreeSans 112 90 0 0 data_in[1]
port 7 nsew signal input
flabel metal2 s 24028 32952 24042 33000 0 FreeSans 112 90 0 0 data_in[2]
port 8 nsew signal input
flabel metal3 s 32920 10763 33000 10793 0 FreeSans 240 0 0 0 data_in[3]
port 9 nsew signal input
flabel metal2 s 23200 32952 23214 33000 0 FreeSans 112 90 0 0 data_in[4]
port 10 nsew signal input
flabel metal2 s 23936 32952 23950 33000 0 FreeSans 112 90 0 0 data_in[5]
port 11 nsew signal input
flabel metal2 s 20532 32952 20546 33000 0 FreeSans 112 90 0 0 data_in[6]
port 12 nsew signal input
flabel metal2 s 21544 32952 21558 33000 0 FreeSans 112 90 0 0 data_in[7]
port 13 nsew signal input
flabel metal2 s 5628 32952 5642 33000 0 FreeSans 112 90 0 0 data_out[0]
port 14 nsew signal output
flabel metal3 s 0 11987 80 12017 0 FreeSans 240 0 0 0 data_out[1]
port 15 nsew signal output
flabel metal2 s 5536 32952 5550 33000 0 FreeSans 112 90 0 0 data_out[2]
port 16 nsew signal output
flabel metal2 s 21084 32952 21098 33000 0 FreeSans 112 90 0 0 data_out[3]
port 17 nsew signal output
flabel metal2 s 13908 0 13922 48 0 FreeSans 112 90 0 0 data_out[4]
port 18 nsew signal output
flabel metal3 s 0 5595 80 5625 0 FreeSans 240 0 0 0 data_out[5]
port 19 nsew signal output
flabel metal2 s 20992 32952 21006 33000 0 FreeSans 112 90 0 0 data_out[6]
port 20 nsew signal output
flabel metal2 s 20900 32952 20914 33000 0 FreeSans 112 90 0 0 data_out[7]
port 21 nsew signal output
flabel metal3 s 0 18515 80 18545 0 FreeSans 240 0 0 0 data_out[8]
port 22 nsew signal output
flabel metal2 s 18692 0 18706 48 0 FreeSans 112 90 0 0 parity_sel
port 23 nsew signal input
flabel metal2 s 19244 32952 19258 33000 0 FreeSans 112 90 0 0 receive
port 24 nsew signal input
flabel metal2 s 14368 32952 14382 33000 0 FreeSans 112 90 0 0 rst
port 25 nsew signal input
flabel metal2 s 16300 0 16314 48 0 FreeSans 112 90 0 0 start_Tx
port 26 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 33000 33000
<< end >>
